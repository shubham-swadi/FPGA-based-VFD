module LUT_method_3(Clk,reset,data_out_3);
    input Clk,reset;
    output reg [11:0] data_out_3;
    reg [20:0] counter; 
    reg [11:0] sine [0:4095];
    integer k;  
    
    initial begin
        k = 0;
sine[0] =34;
sine[1] =34;
sine[2] =34;
sine[3] =34;
sine[4] =33;
sine[5] =33;
sine[6] =33;
sine[7] =33;
sine[8] =33;
sine[9] =32;
sine[10] =32;
sine[11] =32;
sine[12] =32;
sine[13] =32;
sine[14] =31;
sine[15] =31;
sine[16] =31;
sine[17] =31;
sine[18] =31;
sine[19] =31;
sine[20] =30;
sine[21] =30;
sine[22] =30;
sine[23] =30;
sine[24] =30;
sine[25] =29;
sine[26] =29;
sine[27] =29;
sine[28] =29;
sine[29] =29;
sine[30] =29;
sine[31] =28;
sine[32] =28;
sine[33] =28;
sine[34] =28;
sine[35] =28;
sine[36] =27;
sine[37] =27;
sine[38] =27;
sine[39] =27;
sine[40] =27;
sine[41] =27;
sine[42] =26;
sine[43] =26;
sine[44] =26;
sine[45] =26;
sine[46] =26;
sine[47] =26;
sine[48] =25;
sine[49] =25;
sine[50] =25;
sine[51] =25;
sine[52] =25;
sine[53] =25;
sine[54] =24;
sine[55] =24;
sine[56] =24;
sine[57] =24;
sine[58] =24;
sine[59] =24;
sine[60] =23;
sine[61] =23;
sine[62] =23;
sine[63] =23;
sine[64] =23;
sine[65] =23;
sine[66] =22;
sine[67] =22;
sine[68] =22;
sine[69] =22;
sine[70] =22;
sine[71] =22;
sine[72] =21;
sine[73] =21;
sine[74] =21;
sine[75] =21;
sine[76] =21;
sine[77] =21;
sine[78] =21;
sine[79] =20;
sine[80] =20;
sine[81] =20;
sine[82] =20;
sine[83] =20;
sine[84] =20;
sine[85] =19;
sine[86] =19;
sine[87] =19;
sine[88] =19;
sine[89] =19;
sine[90] =19;
sine[91] =19;
sine[92] =18;
sine[93] =18;
sine[94] =18;
sine[95] =18;
sine[96] =18;
sine[97] =18;
sine[98] =18;
sine[99] =17;
sine[100] =17;
sine[101] =17;
sine[102] =17;
sine[103] =17;
sine[104] =17;
sine[105] =17;
sine[106] =16;
sine[107] =16;
sine[108] =16;
sine[109] =16;
sine[110] =16;
sine[111] =16;
sine[112] =16;
sine[113] =15;
sine[114] =15;
sine[115] =15;
sine[116] =15;
sine[117] =15;
sine[118] =15;
sine[119] =15;
sine[120] =15;
sine[121] =14;
sine[122] =14;
sine[123] =14;
sine[124] =14;
sine[125] =14;
sine[126] =14;
sine[127] =14;
sine[128] =14;
sine[129] =13;
sine[130] =13;
sine[131] =13;
sine[132] =13;
sine[133] =13;
sine[134] =13;
sine[135] =13;
sine[136] =13;
sine[137] =12;
sine[138] =12;
sine[139] =12;
sine[140] =12;
sine[141] =12;
sine[142] =12;
sine[143] =12;
sine[144] =12;
sine[145] =11;
sine[146] =11;
sine[147] =11;
sine[148] =11;
sine[149] =11;
sine[150] =11;
sine[151] =11;
sine[152] =11;
sine[153] =11;
sine[154] =10;
sine[155] =10;
sine[156] =10;
sine[157] =10;
sine[158] =10;
sine[159] =10;
sine[160] =10;
sine[161] =10;
sine[162] =10;
sine[163] =9;
sine[164] =9;
sine[165] =9;
sine[166] =9;
sine[167] =9;
sine[168] =9;
sine[169] =9;
sine[170] =9;
sine[171] =9;
sine[172] =9;
sine[173] =8;
sine[174] =8;
sine[175] =8;
sine[176] =8;
sine[177] =8;
sine[178] =8;
sine[179] =8;
sine[180] =8;
sine[181] =8;
sine[182] =8;
sine[183] =7;
sine[184] =7;
sine[185] =7;
sine[186] =7;
sine[187] =7;
sine[188] =7;
sine[189] =7;
sine[190] =7;
sine[191] =7;
sine[192] =7;
sine[193] =7;
sine[194] =6;
sine[195] =6;
sine[196] =6;
sine[197] =6;
sine[198] =6;
sine[199] =6;
sine[200] =6;
sine[201] =6;
sine[202] =6;
sine[203] =6;
sine[204] =6;
sine[205] =6;
sine[206] =5;
sine[207] =5;
sine[208] =5;
sine[209] =5;
sine[210] =5;
sine[211] =5;
sine[212] =5;
sine[213] =5;
sine[214] =5;
sine[215] =5;
sine[216] =5;
sine[217] =5;
sine[218] =5;
sine[219] =4;
sine[220] =4;
sine[221] =4;
sine[222] =4;
sine[223] =4;
sine[224] =4;
sine[225] =4;
sine[226] =4;
sine[227] =4;
sine[228] =4;
sine[229] =4;
sine[230] =4;
sine[231] =4;
sine[232] =4;
sine[233] =3;
sine[234] =3;
sine[235] =3;
sine[236] =3;
sine[237] =3;
sine[238] =3;
sine[239] =3;
sine[240] =3;
sine[241] =3;
sine[242] =3;
sine[243] =3;
sine[244] =3;
sine[245] =3;
sine[246] =3;
sine[247] =3;
sine[248] =3;
sine[249] =3;
sine[250] =2;
sine[251] =2;
sine[252] =2;
sine[253] =2;
sine[254] =2;
sine[255] =2;
sine[256] =2;
sine[257] =2;
sine[258] =2;
sine[259] =2;
sine[260] =2;
sine[261] =2;
sine[262] =2;
sine[263] =2;
sine[264] =2;
sine[265] =2;
sine[266] =2;
sine[267] =2;
sine[268] =2;
sine[269] =2;
sine[270] =2;
sine[271] =1;
sine[272] =1;
sine[273] =1;
sine[274] =1;
sine[275] =1;
sine[276] =1;
sine[277] =1;
sine[278] =1;
sine[279] =1;
sine[280] =1;
sine[281] =1;
sine[282] =1;
sine[283] =1;
sine[284] =1;
sine[285] =1;
sine[286] =1;
sine[287] =1;
sine[288] =1;
sine[289] =1;
sine[290] =1;
sine[291] =1;
sine[292] =1;
sine[293] =1;
sine[294] =1;
sine[295] =1;
sine[296] =1;
sine[297] =1;
sine[298] =1;
sine[299] =1;
sine[300] =1;
sine[301] =0;
sine[302] =0;
sine[303] =0;
sine[304] =0;
sine[305] =0;
sine[306] =0;
sine[307] =0;
sine[308] =0;
sine[309] =0;
sine[310] =0;
sine[311] =0;
sine[312] =0;
sine[313] =0;
sine[314] =0;
sine[315] =0;
sine[316] =0;
sine[317] =0;
sine[318] =0;
sine[319] =0;
sine[320] =0;
sine[321] =0;
sine[322] =0;
sine[323] =0;
sine[324] =0;
sine[325] =0;
sine[326] =0;
sine[327] =0;
sine[328] =0;
sine[329] =0;
sine[330] =0;
sine[331] =0;
sine[332] =0;
sine[333] =0;
sine[334] =0;
sine[335] =0;
sine[336] =0;
sine[337] =0;
sine[338] =0;
sine[339] =0;
sine[340] =0;
sine[341] =0;
sine[342] =0;
sine[343] =0;
sine[344] =0;
sine[345] =0;
sine[346] =0;
sine[347] =0;
sine[348] =0;
sine[349] =0;
sine[350] =0;
sine[351] =0;
sine[352] =0;
sine[353] =0;
sine[354] =0;
sine[355] =0;
sine[356] =0;
sine[357] =0;
sine[358] =0;
sine[359] =0;
sine[360] =0;
sine[361] =0;
sine[362] =0;
sine[363] =0;
sine[364] =0;
sine[365] =0;
sine[366] =0;
sine[367] =0;
sine[368] =0;
sine[369] =0;
sine[370] =0;
sine[371] =0;
sine[372] =0;
sine[373] =0;
sine[374] =0;
sine[375] =0;
sine[376] =0;
sine[377] =0;
sine[378] =0;
sine[379] =0;
sine[380] =0;
sine[381] =0;
sine[382] =1;
sine[383] =1;
sine[384] =1;
sine[385] =1;
sine[386] =1;
sine[387] =1;
sine[388] =1;
sine[389] =1;
sine[390] =1;
sine[391] =1;
sine[392] =1;
sine[393] =1;
sine[394] =1;
sine[395] =1;
sine[396] =1;
sine[397] =1;
sine[398] =1;
sine[399] =1;
sine[400] =1;
sine[401] =1;
sine[402] =1;
sine[403] =1;
sine[404] =1;
sine[405] =1;
sine[406] =1;
sine[407] =1;
sine[408] =1;
sine[409] =1;
sine[410] =1;
sine[411] =1;
sine[412] =2;
sine[413] =2;
sine[414] =2;
sine[415] =2;
sine[416] =2;
sine[417] =2;
sine[418] =2;
sine[419] =2;
sine[420] =2;
sine[421] =2;
sine[422] =2;
sine[423] =2;
sine[424] =2;
sine[425] =2;
sine[426] =2;
sine[427] =2;
sine[428] =2;
sine[429] =2;
sine[430] =2;
sine[431] =2;
sine[432] =2;
sine[433] =3;
sine[434] =3;
sine[435] =3;
sine[436] =3;
sine[437] =3;
sine[438] =3;
sine[439] =3;
sine[440] =3;
sine[441] =3;
sine[442] =3;
sine[443] =3;
sine[444] =3;
sine[445] =3;
sine[446] =3;
sine[447] =3;
sine[448] =3;
sine[449] =3;
sine[450] =4;
sine[451] =4;
sine[452] =4;
sine[453] =4;
sine[454] =4;
sine[455] =4;
sine[456] =4;
sine[457] =4;
sine[458] =4;
sine[459] =4;
sine[460] =4;
sine[461] =4;
sine[462] =4;
sine[463] =4;
sine[464] =5;
sine[465] =5;
sine[466] =5;
sine[467] =5;
sine[468] =5;
sine[469] =5;
sine[470] =5;
sine[471] =5;
sine[472] =5;
sine[473] =5;
sine[474] =5;
sine[475] =5;
sine[476] =5;
sine[477] =6;
sine[478] =6;
sine[479] =6;
sine[480] =6;
sine[481] =6;
sine[482] =6;
sine[483] =6;
sine[484] =6;
sine[485] =6;
sine[486] =6;
sine[487] =6;
sine[488] =6;
sine[489] =7;
sine[490] =7;
sine[491] =7;
sine[492] =7;
sine[493] =7;
sine[494] =7;
sine[495] =7;
sine[496] =7;
sine[497] =7;
sine[498] =7;
sine[499] =7;
sine[500] =8;
sine[501] =8;
sine[502] =8;
sine[503] =8;
sine[504] =8;
sine[505] =8;
sine[506] =8;
sine[507] =8;
sine[508] =8;
sine[509] =8;
sine[510] =9;
sine[511] =9;
sine[512] =9;
sine[513] =9;
sine[514] =9;
sine[515] =9;
sine[516] =9;
sine[517] =9;
sine[518] =9;
sine[519] =9;
sine[520] =10;
sine[521] =10;
sine[522] =10;
sine[523] =10;
sine[524] =10;
sine[525] =10;
sine[526] =10;
sine[527] =10;
sine[528] =10;
sine[529] =11;
sine[530] =11;
sine[531] =11;
sine[532] =11;
sine[533] =11;
sine[534] =11;
sine[535] =11;
sine[536] =11;
sine[537] =11;
sine[538] =12;
sine[539] =12;
sine[540] =12;
sine[541] =12;
sine[542] =12;
sine[543] =12;
sine[544] =12;
sine[545] =12;
sine[546] =13;
sine[547] =13;
sine[548] =13;
sine[549] =13;
sine[550] =13;
sine[551] =13;
sine[552] =13;
sine[553] =13;
sine[554] =14;
sine[555] =14;
sine[556] =14;
sine[557] =14;
sine[558] =14;
sine[559] =14;
sine[560] =14;
sine[561] =14;
sine[562] =15;
sine[563] =15;
sine[564] =15;
sine[565] =15;
sine[566] =15;
sine[567] =15;
sine[568] =15;
sine[569] =15;
sine[570] =16;
sine[571] =16;
sine[572] =16;
sine[573] =16;
sine[574] =16;
sine[575] =16;
sine[576] =16;
sine[577] =17;
sine[578] =17;
sine[579] =17;
sine[580] =17;
sine[581] =17;
sine[582] =17;
sine[583] =17;
sine[584] =18;
sine[585] =18;
sine[586] =18;
sine[587] =18;
sine[588] =18;
sine[589] =18;
sine[590] =18;
sine[591] =19;
sine[592] =19;
sine[593] =19;
sine[594] =19;
sine[595] =19;
sine[596] =19;
sine[597] =19;
sine[598] =20;
sine[599] =20;
sine[600] =20;
sine[601] =20;
sine[602] =20;
sine[603] =20;
sine[604] =21;
sine[605] =21;
sine[606] =21;
sine[607] =21;
sine[608] =21;
sine[609] =21;
sine[610] =21;
sine[611] =22;
sine[612] =22;
sine[613] =22;
sine[614] =22;
sine[615] =22;
sine[616] =22;
sine[617] =23;
sine[618] =23;
sine[619] =23;
sine[620] =23;
sine[621] =23;
sine[622] =23;
sine[623] =24;
sine[624] =24;
sine[625] =24;
sine[626] =24;
sine[627] =24;
sine[628] =24;
sine[629] =25;
sine[630] =25;
sine[631] =25;
sine[632] =25;
sine[633] =25;
sine[634] =25;
sine[635] =26;
sine[636] =26;
sine[637] =26;
sine[638] =26;
sine[639] =26;
sine[640] =26;
sine[641] =27;
sine[642] =27;
sine[643] =27;
sine[644] =27;
sine[645] =27;
sine[646] =27;
sine[647] =28;
sine[648] =28;
sine[649] =28;
sine[650] =28;
sine[651] =28;
sine[652] =29;
sine[653] =29;
sine[654] =29;
sine[655] =29;
sine[656] =29;
sine[657] =29;
sine[658] =30;
sine[659] =30;
sine[660] =30;
sine[661] =30;
sine[662] =30;
sine[663] =31;
sine[664] =31;
sine[665] =31;
sine[666] =31;
sine[667] =31;
sine[668] =31;
sine[669] =32;
sine[670] =32;
sine[671] =32;
sine[672] =32;
sine[673] =32;
sine[674] =33;
sine[675] =33;
sine[676] =33;
sine[677] =33;
sine[678] =33;
sine[679] =34;
sine[680] =34;
sine[681] =34;
sine[682] =34;
sine[683] =34;
sine[684] =35;
sine[685] =35;
sine[686] =35;
sine[687] =35;
sine[688] =35;
sine[689] =36;
sine[690] =36;
sine[691] =36;
sine[692] =36;
sine[693] =36;
sine[694] =37;
sine[695] =37;
sine[696] =37;
sine[697] =37;
sine[698] =37;
sine[699] =38;
sine[700] =38;
sine[701] =38;
sine[702] =38;
sine[703] =38;
sine[704] =39;
sine[705] =39;
sine[706] =39;
sine[707] =39;
sine[708] =39;
sine[709] =40;
sine[710] =40;
sine[711] =40;
sine[712] =40;
sine[713] =40;
sine[714] =41;
sine[715] =41;
sine[716] =41;
sine[717] =41;
sine[718] =42;
sine[719] =42;
sine[720] =42;
sine[721] =42;
sine[722] =42;
sine[723] =43;
sine[724] =43;
sine[725] =43;
sine[726] =43;
sine[727] =43;
sine[728] =44;
sine[729] =44;
sine[730] =44;
sine[731] =44;
sine[732] =45;
sine[733] =45;
sine[734] =45;
sine[735] =45;
sine[736] =45;
sine[737] =46;
sine[738] =46;
sine[739] =46;
sine[740] =46;
sine[741] =47;
sine[742] =47;
sine[743] =47;
sine[744] =47;
sine[745] =48;
sine[746] =48;
sine[747] =48;
sine[748] =48;
sine[749] =48;
sine[750] =49;
sine[751] =49;
sine[752] =49;
sine[753] =49;
sine[754] =50;
sine[755] =50;
sine[756] =50;
sine[757] =50;
sine[758] =51;
sine[759] =51;
sine[760] =51;
sine[761] =51;
sine[762] =51;
sine[763] =52;
sine[764] =52;
sine[765] =52;
sine[766] =52;
sine[767] =53;
sine[768] =53;
sine[769] =53;
sine[770] =53;
sine[771] =54;
sine[772] =54;
sine[773] =54;
sine[774] =54;
sine[775] =55;
sine[776] =55;
sine[777] =55;
sine[778] =55;
sine[779] =56;
sine[780] =56;
sine[781] =56;
sine[782] =56;
sine[783] =57;
sine[784] =57;
sine[785] =57;
sine[786] =57;
sine[787] =57;
sine[788] =58;
sine[789] =58;
sine[790] =58;
sine[791] =58;
sine[792] =59;
sine[793] =59;
sine[794] =59;
sine[795] =59;
sine[796] =60;
sine[797] =60;
sine[798] =60;
sine[799] =61;
sine[800] =61;
sine[801] =61;
sine[802] =61;
sine[803] =62;
sine[804] =62;
sine[805] =62;
sine[806] =62;
sine[807] =63;
sine[808] =63;
sine[809] =63;
sine[810] =63;
sine[811] =64;
sine[812] =64;
sine[813] =64;
sine[814] =64;
sine[815] =65;
sine[816] =65;
sine[817] =65;
sine[818] =65;
sine[819] =66;
sine[820] =66;
sine[821] =66;
sine[822] =66;
sine[823] =67;
sine[824] =67;
sine[825] =67;
sine[826] =68;
sine[827] =68;
sine[828] =68;
sine[829] =68;
sine[830] =69;
sine[831] =69;
sine[832] =69;
sine[833] =69;
sine[834] =70;
sine[835] =70;
sine[836] =70;
sine[837] =70;
sine[838] =71;
sine[839] =71;
sine[840] =71;
sine[841] =72;
sine[842] =72;
sine[843] =72;
sine[844] =72;
sine[845] =73;
sine[846] =73;
sine[847] =73;
sine[848] =73;
sine[849] =74;
sine[850] =74;
sine[851] =74;
sine[852] =75;
sine[853] =75;
sine[854] =75;
sine[855] =75;
sine[856] =76;
sine[857] =76;
sine[858] =76;
sine[859] =77;
sine[860] =77;
sine[861] =77;
sine[862] =77;
sine[863] =78;
sine[864] =78;
sine[865] =78;
sine[866] =78;
sine[867] =79;
sine[868] =79;
sine[869] =79;
sine[870] =80;
sine[871] =80;
sine[872] =80;
sine[873] =80;
sine[874] =81;
sine[875] =81;
sine[876] =81;
sine[877] =82;
sine[878] =82;
sine[879] =82;
sine[880] =82;
sine[881] =83;
sine[882] =83;
sine[883] =83;
sine[884] =84;
sine[885] =84;
sine[886] =84;
sine[887] =84;
sine[888] =85;
sine[889] =85;
sine[890] =85;
sine[891] =86;
sine[892] =86;
sine[893] =86;
sine[894] =87;
sine[895] =87;
sine[896] =87;
sine[897] =87;
sine[898] =88;
sine[899] =88;
sine[900] =88;
sine[901] =89;
sine[902] =89;
sine[903] =89;
sine[904] =90;
sine[905] =90;
sine[906] =90;
sine[907] =90;
sine[908] =91;
sine[909] =91;
sine[910] =91;
sine[911] =92;
sine[912] =92;
sine[913] =92;
sine[914] =93;
sine[915] =93;
sine[916] =93;
sine[917] =93;
sine[918] =94;
sine[919] =94;
sine[920] =94;
sine[921] =95;
sine[922] =95;
sine[923] =95;
sine[924] =96;
sine[925] =96;
sine[926] =96;
sine[927] =96;
sine[928] =97;
sine[929] =97;
sine[930] =97;
sine[931] =98;
sine[932] =98;
sine[933] =98;
sine[934] =99;
sine[935] =99;
sine[936] =99;
sine[937] =100;
sine[938] =100;
sine[939] =100;
sine[940] =100;
sine[941] =101;
sine[942] =101;
sine[943] =101;
sine[944] =102;
sine[945] =102;
sine[946] =102;
sine[947] =103;
sine[948] =103;
sine[949] =103;
sine[950] =104;
sine[951] =104;
sine[952] =104;
sine[953] =105;
sine[954] =105;
sine[955] =105;
sine[956] =106;
sine[957] =106;
sine[958] =106;
sine[959] =106;
sine[960] =107;
sine[961] =107;
sine[962] =107;
sine[963] =108;
sine[964] =108;
sine[965] =108;
sine[966] =109;
sine[967] =109;
sine[968] =109;
sine[969] =110;
sine[970] =110;
sine[971] =110;
sine[972] =111;
sine[973] =111;
sine[974] =111;
sine[975] =112;
sine[976] =112;
sine[977] =112;
sine[978] =113;
sine[979] =113;
sine[980] =113;
sine[981] =114;
sine[982] =114;
sine[983] =114;
sine[984] =115;
sine[985] =115;
sine[986] =115;
sine[987] =116;
sine[988] =116;
sine[989] =116;
sine[990] =116;
sine[991] =117;
sine[992] =117;
sine[993] =117;
sine[994] =118;
sine[995] =118;
sine[996] =118;
sine[997] =119;
sine[998] =119;
sine[999] =119;
sine[1000] =120;
sine[1001] =120;
sine[1002] =120;
sine[1003] =121;
sine[1004] =121;
sine[1005] =121;
sine[1006] =122;
sine[1007] =122;
sine[1008] =122;
sine[1009] =123;
sine[1010] =123;
sine[1011] =123;
sine[1012] =124;
sine[1013] =124;
sine[1014] =124;
sine[1015] =125;
sine[1016] =125;
sine[1017] =125;
sine[1018] =126;
sine[1019] =126;
sine[1020] =127;
sine[1021] =127;
sine[1022] =127;
sine[1023] =128;
sine[1024] =128;
sine[1025] =128;
sine[1026] =129;
sine[1027] =129;
sine[1028] =129;
sine[1029] =130;
sine[1030] =130;
sine[1031] =130;
sine[1032] =131;
sine[1033] =131;
sine[1034] =131;
sine[1035] =132;
sine[1036] =132;
sine[1037] =132;
sine[1038] =133;
sine[1039] =133;
sine[1040] =133;
sine[1041] =134;
sine[1042] =134;
sine[1043] =134;
sine[1044] =135;
sine[1045] =135;
sine[1046] =135;
sine[1047] =136;
sine[1048] =136;
sine[1049] =136;
sine[1050] =137;
sine[1051] =137;
sine[1052] =137;
sine[1053] =138;
sine[1054] =138;
sine[1055] =139;
sine[1056] =139;
sine[1057] =139;
sine[1058] =140;
sine[1059] =140;
sine[1060] =140;
sine[1061] =141;
sine[1062] =141;
sine[1063] =141;
sine[1064] =142;
sine[1065] =142;
sine[1066] =142;
sine[1067] =143;
sine[1068] =143;
sine[1069] =143;
sine[1070] =144;
sine[1071] =144;
sine[1072] =144;
sine[1073] =145;
sine[1074] =145;
sine[1075] =146;
sine[1076] =146;
sine[1077] =146;
sine[1078] =147;
sine[1079] =147;
sine[1080] =147;
sine[1081] =148;
sine[1082] =148;
sine[1083] =148;
sine[1084] =149;
sine[1085] =149;
sine[1086] =149;
sine[1087] =150;
sine[1088] =150;
sine[1089] =151;
sine[1090] =151;
sine[1091] =151;
sine[1092] =152;
sine[1093] =152;
sine[1094] =152;
sine[1095] =153;
sine[1096] =153;
sine[1097] =153;
sine[1098] =154;
sine[1099] =154;
sine[1100] =154;
sine[1101] =155;
sine[1102] =155;
sine[1103] =156;
sine[1104] =156;
sine[1105] =156;
sine[1106] =157;
sine[1107] =157;
sine[1108] =157;
sine[1109] =158;
sine[1110] =158;
sine[1111] =158;
sine[1112] =159;
sine[1113] =159;
sine[1114] =160;
sine[1115] =160;
sine[1116] =160;
sine[1117] =161;
sine[1118] =161;
sine[1119] =161;
sine[1120] =162;
sine[1121] =162;
sine[1122] =162;
sine[1123] =163;
sine[1124] =163;
sine[1125] =164;
sine[1126] =164;
sine[1127] =164;
sine[1128] =165;
sine[1129] =165;
sine[1130] =165;
sine[1131] =166;
sine[1132] =166;
sine[1133] =166;
sine[1134] =167;
sine[1135] =167;
sine[1136] =168;
sine[1137] =168;
sine[1138] =168;
sine[1139] =169;
sine[1140] =169;
sine[1141] =169;
sine[1142] =170;
sine[1143] =170;
sine[1144] =171;
sine[1145] =171;
sine[1146] =171;
sine[1147] =172;
sine[1148] =172;
sine[1149] =172;
sine[1150] =173;
sine[1151] =173;
sine[1152] =173;
sine[1153] =174;
sine[1154] =174;
sine[1155] =175;
sine[1156] =175;
sine[1157] =175;
sine[1158] =176;
sine[1159] =176;
sine[1160] =176;
sine[1161] =177;
sine[1162] =177;
sine[1163] =178;
sine[1164] =178;
sine[1165] =178;
sine[1166] =179;
sine[1167] =179;
sine[1168] =179;
sine[1169] =180;
sine[1170] =180;
sine[1171] =181;
sine[1172] =181;
sine[1173] =181;
sine[1174] =182;
sine[1175] =182;
sine[1176] =182;
sine[1177] =183;
sine[1178] =183;
sine[1179] =184;
sine[1180] =184;
sine[1181] =184;
sine[1182] =185;
sine[1183] =185;
sine[1184] =185;
sine[1185] =186;
sine[1186] =186;
sine[1187] =187;
sine[1188] =187;
sine[1189] =187;
sine[1190] =188;
sine[1191] =188;
sine[1192] =188;
sine[1193] =189;
sine[1194] =189;
sine[1195] =190;
sine[1196] =190;
sine[1197] =190;
sine[1198] =191;
sine[1199] =191;
sine[1200] =192;
sine[1201] =192;
sine[1202] =192;
sine[1203] =193;
sine[1204] =193;
sine[1205] =193;
sine[1206] =194;
sine[1207] =194;
sine[1208] =195;
sine[1209] =195;
sine[1210] =195;
sine[1211] =196;
sine[1212] =196;
sine[1213] =196;
sine[1214] =197;
sine[1215] =197;
sine[1216] =198;
sine[1217] =198;
sine[1218] =198;
sine[1219] =199;
sine[1220] =199;
sine[1221] =200;
sine[1222] =200;
sine[1223] =200;
sine[1224] =201;
sine[1225] =201;
sine[1226] =201;
sine[1227] =202;
sine[1228] =202;
sine[1229] =203;
sine[1230] =203;
sine[1231] =203;
sine[1232] =204;
sine[1233] =204;
sine[1234] =205;
sine[1235] =205;
sine[1236] =205;
sine[1237] =206;
sine[1238] =206;
sine[1239] =206;
sine[1240] =207;
sine[1241] =207;
sine[1242] =208;
sine[1243] =208;
sine[1244] =208;
sine[1245] =209;
sine[1246] =209;
sine[1247] =210;
sine[1248] =210;
sine[1249] =210;
sine[1250] =211;
sine[1251] =211;
sine[1252] =211;
sine[1253] =212;
sine[1254] =212;
sine[1255] =213;
sine[1256] =213;
sine[1257] =213;
sine[1258] =214;
sine[1259] =214;
sine[1260] =215;
sine[1261] =215;
sine[1262] =215;
sine[1263] =216;
sine[1264] =216;
sine[1265] =216;
sine[1266] =217;
sine[1267] =217;
sine[1268] =218;
sine[1269] =218;
sine[1270] =218;
sine[1271] =219;
sine[1272] =219;
sine[1273] =220;
sine[1274] =220;
sine[1275] =220;
sine[1276] =221;
sine[1277] =221;
sine[1278] =222;
sine[1279] =222;
sine[1280] =222;
sine[1281] =223;
sine[1282] =223;
sine[1283] =223;
sine[1284] =224;
sine[1285] =224;
sine[1286] =225;
sine[1287] =225;
sine[1288] =225;
sine[1289] =226;
sine[1290] =226;
sine[1291] =227;
sine[1292] =227;
sine[1293] =227;
sine[1294] =228;
sine[1295] =228;
sine[1296] =229;
sine[1297] =229;
sine[1298] =229;
sine[1299] =230;
sine[1300] =230;
sine[1301] =230;
sine[1302] =231;
sine[1303] =231;
sine[1304] =232;
sine[1305] =232;
sine[1306] =232;
sine[1307] =233;
sine[1308] =233;
sine[1309] =234;
sine[1310] =234;
sine[1311] =234;
sine[1312] =235;
sine[1313] =235;
sine[1314] =236;
sine[1315] =236;
sine[1316] =236;
sine[1317] =237;
sine[1318] =237;
sine[1319] =237;
sine[1320] =238;
sine[1321] =238;
sine[1322] =239;
sine[1323] =239;
sine[1324] =239;
sine[1325] =240;
sine[1326] =240;
sine[1327] =241;
sine[1328] =241;
sine[1329] =241;
sine[1330] =242;
sine[1331] =242;
sine[1332] =243;
sine[1333] =243;
sine[1334] =243;
sine[1335] =244;
sine[1336] =244;
sine[1337] =245;
sine[1338] =245;
sine[1339] =245;
sine[1340] =246;
sine[1341] =246;
sine[1342] =246;
sine[1343] =247;
sine[1344] =247;
sine[1345] =248;
sine[1346] =248;
sine[1347] =248;
sine[1348] =249;
sine[1349] =249;
sine[1350] =250;
sine[1351] =250;
sine[1352] =250;
sine[1353] =251;
sine[1354] =251;
sine[1355] =252;
sine[1356] =252;
sine[1357] =252;
sine[1358] =253;
sine[1359] =253;
sine[1360] =254;
sine[1361] =254;
sine[1362] =254;
sine[1363] =255;
sine[1364] =255;
sine[1365] =256;
sine[1366] =256;
sine[1367] =256;
sine[1368] =257;
sine[1369] =257;
sine[1370] =257;
sine[1371] =258;
sine[1372] =258;
sine[1373] =259;
sine[1374] =259;
sine[1375] =259;
sine[1376] =260;
sine[1377] =260;
sine[1378] =261;
sine[1379] =261;
sine[1380] =261;
sine[1381] =262;
sine[1382] =262;
sine[1383] =263;
sine[1384] =263;
sine[1385] =263;
sine[1386] =264;
sine[1387] =264;
sine[1388] =265;
sine[1389] =265;
sine[1390] =265;
sine[1391] =266;
sine[1392] =266;
sine[1393] =266;
sine[1394] =267;
sine[1395] =267;
sine[1396] =268;
sine[1397] =268;
sine[1398] =268;
sine[1399] =269;
sine[1400] =269;
sine[1401] =270;
sine[1402] =270;
sine[1403] =270;
sine[1404] =271;
sine[1405] =271;
sine[1406] =272;
sine[1407] =272;
sine[1408] =272;
sine[1409] =273;
sine[1410] =273;
sine[1411] =274;
sine[1412] =274;
sine[1413] =274;
sine[1414] =275;
sine[1415] =275;
sine[1416] =275;
sine[1417] =276;
sine[1418] =276;
sine[1419] =277;
sine[1420] =277;
sine[1421] =277;
sine[1422] =278;
sine[1423] =278;
sine[1424] =279;
sine[1425] =279;
sine[1426] =279;
sine[1427] =280;
sine[1428] =280;
sine[1429] =281;
sine[1430] =281;
sine[1431] =281;
sine[1432] =282;
sine[1433] =282;
sine[1434] =282;
sine[1435] =283;
sine[1436] =283;
sine[1437] =284;
sine[1438] =284;
sine[1439] =284;
sine[1440] =285;
sine[1441] =285;
sine[1442] =286;
sine[1443] =286;
sine[1444] =286;
sine[1445] =287;
sine[1446] =287;
sine[1447] =288;
sine[1448] =288;
sine[1449] =288;
sine[1450] =289;
sine[1451] =289;
sine[1452] =289;
sine[1453] =290;
sine[1454] =290;
sine[1455] =291;
sine[1456] =291;
sine[1457] =291;
sine[1458] =292;
sine[1459] =292;
sine[1460] =293;
sine[1461] =293;
sine[1462] =293;
sine[1463] =294;
sine[1464] =294;
sine[1465] =295;
sine[1466] =295;
sine[1467] =295;
sine[1468] =296;
sine[1469] =296;
sine[1470] =296;
sine[1471] =297;
sine[1472] =297;
sine[1473] =298;
sine[1474] =298;
sine[1475] =298;
sine[1476] =299;
sine[1477] =299;
sine[1478] =300;
sine[1479] =300;
sine[1480] =300;
sine[1481] =301;
sine[1482] =301;
sine[1483] =301;
sine[1484] =302;
sine[1485] =302;
sine[1486] =303;
sine[1487] =303;
sine[1488] =303;
sine[1489] =304;
sine[1490] =304;
sine[1491] =305;
sine[1492] =305;
sine[1493] =305;
sine[1494] =306;
sine[1495] =306;
sine[1496] =306;
sine[1497] =307;
sine[1498] =307;
sine[1499] =308;
sine[1500] =308;
sine[1501] =308;
sine[1502] =309;
sine[1503] =309;
sine[1504] =310;
sine[1505] =310;
sine[1506] =310;
sine[1507] =311;
sine[1508] =311;
sine[1509] =311;
sine[1510] =312;
sine[1511] =312;
sine[1512] =313;
sine[1513] =313;
sine[1514] =313;
sine[1515] =314;
sine[1516] =314;
sine[1517] =315;
sine[1518] =315;
sine[1519] =315;
sine[1520] =316;
sine[1521] =316;
sine[1522] =316;
sine[1523] =317;
sine[1524] =317;
sine[1525] =318;
sine[1526] =318;
sine[1527] =318;
sine[1528] =319;
sine[1529] =319;
sine[1530] =319;
sine[1531] =320;
sine[1532] =320;
sine[1533] =321;
sine[1534] =321;
sine[1535] =321;
sine[1536] =322;
sine[1537] =322;
sine[1538] =323;
sine[1539] =323;
sine[1540] =323;
sine[1541] =324;
sine[1542] =324;
sine[1543] =324;
sine[1544] =325;
sine[1545] =325;
sine[1546] =326;
sine[1547] =326;
sine[1548] =326;
sine[1549] =327;
sine[1550] =327;
sine[1551] =327;
sine[1552] =328;
sine[1553] =328;
sine[1554] =329;
sine[1555] =329;
sine[1556] =329;
sine[1557] =330;
sine[1558] =330;
sine[1559] =330;
sine[1560] =331;
sine[1561] =331;
sine[1562] =332;
sine[1563] =332;
sine[1564] =332;
sine[1565] =333;
sine[1566] =333;
sine[1567] =333;
sine[1568] =334;
sine[1569] =334;
sine[1570] =335;
sine[1571] =335;
sine[1572] =335;
sine[1573] =336;
sine[1574] =336;
sine[1575] =336;
sine[1576] =337;
sine[1577] =337;
sine[1578] =338;
sine[1579] =338;
sine[1580] =338;
sine[1581] =339;
sine[1582] =339;
sine[1583] =339;
sine[1584] =340;
sine[1585] =340;
sine[1586] =340;
sine[1587] =341;
sine[1588] =341;
sine[1589] =342;
sine[1590] =342;
sine[1591] =342;
sine[1592] =343;
sine[1593] =343;
sine[1594] =343;
sine[1595] =344;
sine[1596] =344;
sine[1597] =345;
sine[1598] =345;
sine[1599] =345;
sine[1600] =346;
sine[1601] =346;
sine[1602] =346;
sine[1603] =347;
sine[1604] =347;
sine[1605] =347;
sine[1606] =348;
sine[1607] =348;
sine[1608] =349;
sine[1609] =349;
sine[1610] =349;
sine[1611] =350;
sine[1612] =350;
sine[1613] =350;
sine[1614] =351;
sine[1615] =351;
sine[1616] =351;
sine[1617] =352;
sine[1618] =352;
sine[1619] =353;
sine[1620] =353;
sine[1621] =353;
sine[1622] =354;
sine[1623] =354;
sine[1624] =354;
sine[1625] =355;
sine[1626] =355;
sine[1627] =355;
sine[1628] =356;
sine[1629] =356;
sine[1630] =357;
sine[1631] =357;
sine[1632] =357;
sine[1633] =358;
sine[1634] =358;
sine[1635] =358;
sine[1636] =359;
sine[1637] =359;
sine[1638] =359;
sine[1639] =360;
sine[1640] =360;
sine[1641] =360;
sine[1642] =361;
sine[1643] =361;
sine[1644] =362;
sine[1645] =362;
sine[1646] =362;
sine[1647] =363;
sine[1648] =363;
sine[1649] =363;
sine[1650] =364;
sine[1651] =364;
sine[1652] =364;
sine[1653] =365;
sine[1654] =365;
sine[1655] =365;
sine[1656] =366;
sine[1657] =366;
sine[1658] =367;
sine[1659] =367;
sine[1660] =367;
sine[1661] =368;
sine[1662] =368;
sine[1663] =368;
sine[1664] =369;
sine[1665] =369;
sine[1666] =369;
sine[1667] =370;
sine[1668] =370;
sine[1669] =370;
sine[1670] =371;
sine[1671] =371;
sine[1672] =371;
sine[1673] =372;
sine[1674] =372;
sine[1675] =372;
sine[1676] =373;
sine[1677] =373;
sine[1678] =374;
sine[1679] =374;
sine[1680] =374;
sine[1681] =375;
sine[1682] =375;
sine[1683] =375;
sine[1684] =376;
sine[1685] =376;
sine[1686] =376;
sine[1687] =377;
sine[1688] =377;
sine[1689] =377;
sine[1690] =378;
sine[1691] =378;
sine[1692] =378;
sine[1693] =379;
sine[1694] =379;
sine[1695] =379;
sine[1696] =380;
sine[1697] =380;
sine[1698] =380;
sine[1699] =381;
sine[1700] =381;
sine[1701] =381;
sine[1702] =382;
sine[1703] =382;
sine[1704] =382;
sine[1705] =383;
sine[1706] =383;
sine[1707] =383;
sine[1708] =384;
sine[1709] =384;
sine[1710] =384;
sine[1711] =385;
sine[1712] =385;
sine[1713] =386;
sine[1714] =386;
sine[1715] =386;
sine[1716] =387;
sine[1717] =387;
sine[1718] =387;
sine[1719] =388;
sine[1720] =388;
sine[1721] =388;
sine[1722] =389;
sine[1723] =389;
sine[1724] =389;
sine[1725] =390;
sine[1726] =390;
sine[1727] =390;
sine[1728] =391;
sine[1729] =391;
sine[1730] =391;
sine[1731] =392;
sine[1732] =392;
sine[1733] =392;
sine[1734] =393;
sine[1735] =393;
sine[1736] =393;
sine[1737] =394;
sine[1738] =394;
sine[1739] =394;
sine[1740] =395;
sine[1741] =395;
sine[1742] =395;
sine[1743] =395;
sine[1744] =396;
sine[1745] =396;
sine[1746] =396;
sine[1747] =397;
sine[1748] =397;
sine[1749] =397;
sine[1750] =398;
sine[1751] =398;
sine[1752] =398;
sine[1753] =399;
sine[1754] =399;
sine[1755] =399;
sine[1756] =400;
sine[1757] =400;
sine[1758] =400;
sine[1759] =401;
sine[1760] =401;
sine[1761] =401;
sine[1762] =402;
sine[1763] =402;
sine[1764] =402;
sine[1765] =403;
sine[1766] =403;
sine[1767] =403;
sine[1768] =404;
sine[1769] =404;
sine[1770] =404;
sine[1771] =405;
sine[1772] =405;
sine[1773] =405;
sine[1774] =405;
sine[1775] =406;
sine[1776] =406;
sine[1777] =406;
sine[1778] =407;
sine[1779] =407;
sine[1780] =407;
sine[1781] =408;
sine[1782] =408;
sine[1783] =408;
sine[1784] =409;
sine[1785] =409;
sine[1786] =409;
sine[1787] =410;
sine[1788] =410;
sine[1789] =410;
sine[1790] =411;
sine[1791] =411;
sine[1792] =411;
sine[1793] =411;
sine[1794] =412;
sine[1795] =412;
sine[1796] =412;
sine[1797] =413;
sine[1798] =413;
sine[1799] =413;
sine[1800] =414;
sine[1801] =414;
sine[1802] =414;
sine[1803] =415;
sine[1804] =415;
sine[1805] =415;
sine[1806] =415;
sine[1807] =416;
sine[1808] =416;
sine[1809] =416;
sine[1810] =417;
sine[1811] =417;
sine[1812] =417;
sine[1813] =418;
sine[1814] =418;
sine[1815] =418;
sine[1816] =418;
sine[1817] =419;
sine[1818] =419;
sine[1819] =419;
sine[1820] =420;
sine[1821] =420;
sine[1822] =420;
sine[1823] =421;
sine[1824] =421;
sine[1825] =421;
sine[1826] =421;
sine[1827] =422;
sine[1828] =422;
sine[1829] =422;
sine[1830] =423;
sine[1831] =423;
sine[1832] =423;
sine[1833] =424;
sine[1834] =424;
sine[1835] =424;
sine[1836] =424;
sine[1837] =425;
sine[1838] =425;
sine[1839] =425;
sine[1840] =426;
sine[1841] =426;
sine[1842] =426;
sine[1843] =427;
sine[1844] =427;
sine[1845] =427;
sine[1846] =427;
sine[1847] =428;
sine[1848] =428;
sine[1849] =428;
sine[1850] =429;
sine[1851] =429;
sine[1852] =429;
sine[1853] =429;
sine[1854] =430;
sine[1855] =430;
sine[1856] =430;
sine[1857] =431;
sine[1858] =431;
sine[1859] =431;
sine[1860] =431;
sine[1861] =432;
sine[1862] =432;
sine[1863] =432;
sine[1864] =433;
sine[1865] =433;
sine[1866] =433;
sine[1867] =433;
sine[1868] =434;
sine[1869] =434;
sine[1870] =434;
sine[1871] =434;
sine[1872] =435;
sine[1873] =435;
sine[1874] =435;
sine[1875] =436;
sine[1876] =436;
sine[1877] =436;
sine[1878] =436;
sine[1879] =437;
sine[1880] =437;
sine[1881] =437;
sine[1882] =438;
sine[1883] =438;
sine[1884] =438;
sine[1885] =438;
sine[1886] =439;
sine[1887] =439;
sine[1888] =439;
sine[1889] =439;
sine[1890] =440;
sine[1891] =440;
sine[1892] =440;
sine[1893] =441;
sine[1894] =441;
sine[1895] =441;
sine[1896] =441;
sine[1897] =442;
sine[1898] =442;
sine[1899] =442;
sine[1900] =442;
sine[1901] =443;
sine[1902] =443;
sine[1903] =443;
sine[1904] =443;
sine[1905] =444;
sine[1906] =444;
sine[1907] =444;
sine[1908] =445;
sine[1909] =445;
sine[1910] =445;
sine[1911] =445;
sine[1912] =446;
sine[1913] =446;
sine[1914] =446;
sine[1915] =446;
sine[1916] =447;
sine[1917] =447;
sine[1918] =447;
sine[1919] =447;
sine[1920] =448;
sine[1921] =448;
sine[1922] =448;
sine[1923] =448;
sine[1924] =449;
sine[1925] =449;
sine[1926] =449;
sine[1927] =449;
sine[1928] =450;
sine[1929] =450;
sine[1930] =450;
sine[1931] =450;
sine[1932] =451;
sine[1933] =451;
sine[1934] =451;
sine[1935] =452;
sine[1936] =452;
sine[1937] =452;
sine[1938] =452;
sine[1939] =453;
sine[1940] =453;
sine[1941] =453;
sine[1942] =453;
sine[1943] =454;
sine[1944] =454;
sine[1945] =454;
sine[1946] =454;
sine[1947] =454;
sine[1948] =455;
sine[1949] =455;
sine[1950] =455;
sine[1951] =455;
sine[1952] =456;
sine[1953] =456;
sine[1954] =456;
sine[1955] =456;
sine[1956] =457;
sine[1957] =457;
sine[1958] =457;
sine[1959] =457;
sine[1960] =458;
sine[1961] =458;
sine[1962] =458;
sine[1963] =458;
sine[1964] =459;
sine[1965] =459;
sine[1966] =459;
sine[1967] =459;
sine[1968] =460;
sine[1969] =460;
sine[1970] =460;
sine[1971] =460;
sine[1972] =460;
sine[1973] =461;
sine[1974] =461;
sine[1975] =461;
sine[1976] =461;
sine[1977] =462;
sine[1978] =462;
sine[1979] =462;
sine[1980] =462;
sine[1981] =463;
sine[1982] =463;
sine[1983] =463;
sine[1984] =463;
sine[1985] =463;
sine[1986] =464;
sine[1987] =464;
sine[1988] =464;
sine[1989] =464;
sine[1990] =465;
sine[1991] =465;
sine[1992] =465;
sine[1993] =465;
sine[1994] =466;
sine[1995] =466;
sine[1996] =466;
sine[1997] =466;
sine[1998] =466;
sine[1999] =467;
sine[2000] =467;
sine[2001] =467;
sine[2002] =467;
sine[2003] =468;
sine[2004] =468;
sine[2005] =468;
sine[2006] =468;
sine[2007] =468;
sine[2008] =469;
sine[2009] =469;
sine[2010] =469;
sine[2011] =469;
sine[2012] =469;
sine[2013] =470;
sine[2014] =470;
sine[2015] =470;
sine[2016] =470;
sine[2017] =471;
sine[2018] =471;
sine[2019] =471;
sine[2020] =471;
sine[2021] =471;
sine[2022] =472;
sine[2023] =472;
sine[2024] =472;
sine[2025] =472;
sine[2026] =472;
sine[2027] =473;
sine[2028] =473;
sine[2029] =473;
sine[2030] =473;
sine[2031] =473;
sine[2032] =474;
sine[2033] =474;
sine[2034] =474;
sine[2035] =474;
sine[2036] =474;
sine[2037] =475;
sine[2038] =475;
sine[2039] =475;
sine[2040] =475;
sine[2041] =475;
sine[2042] =476;
sine[2043] =476;
sine[2044] =476;
sine[2045] =476;
sine[2046] =476;
sine[2047] =477;
sine[2048] =477;
sine[2049] =477;
sine[2050] =477;
sine[2051] =477;
sine[2052] =478;
sine[2053] =478;
sine[2054] =478;
sine[2055] =478;
sine[2056] =478;
sine[2057] =479;
sine[2058] =479;
sine[2059] =479;
sine[2060] =479;
sine[2061] =479;
sine[2062] =480;
sine[2063] =480;
sine[2064] =480;
sine[2065] =480;
sine[2066] =480;
sine[2067] =480;
sine[2068] =481;
sine[2069] =481;
sine[2070] =481;
sine[2071] =481;
sine[2072] =481;
sine[2073] =482;
sine[2074] =482;
sine[2075] =482;
sine[2076] =482;
sine[2077] =482;
sine[2078] =482;
sine[2079] =483;
sine[2080] =483;
sine[2081] =483;
sine[2082] =483;
sine[2083] =483;
sine[2084] =484;
sine[2085] =484;
sine[2086] =484;
sine[2087] =484;
sine[2088] =484;
sine[2089] =484;
sine[2090] =485;
sine[2091] =485;
sine[2092] =485;
sine[2093] =485;
sine[2094] =485;
sine[2095] =485;
sine[2096] =486;
sine[2097] =486;
sine[2098] =486;
sine[2099] =486;
sine[2100] =486;
sine[2101] =486;
sine[2102] =487;
sine[2103] =487;
sine[2104] =487;
sine[2105] =487;
sine[2106] =487;
sine[2107] =487;
sine[2108] =488;
sine[2109] =488;
sine[2110] =488;
sine[2111] =488;
sine[2112] =488;
sine[2113] =488;
sine[2114] =489;
sine[2115] =489;
sine[2116] =489;
sine[2117] =489;
sine[2118] =489;
sine[2119] =489;
sine[2120] =490;
sine[2121] =490;
sine[2122] =490;
sine[2123] =490;
sine[2124] =490;
sine[2125] =490;
sine[2126] =490;
sine[2127] =491;
sine[2128] =491;
sine[2129] =491;
sine[2130] =491;
sine[2131] =491;
sine[2132] =491;
sine[2133] =492;
sine[2134] =492;
sine[2135] =492;
sine[2136] =492;
sine[2137] =492;
sine[2138] =492;
sine[2139] =492;
sine[2140] =493;
sine[2141] =493;
sine[2142] =493;
sine[2143] =493;
sine[2144] =493;
sine[2145] =493;
sine[2146] =493;
sine[2147] =494;
sine[2148] =494;
sine[2149] =494;
sine[2150] =494;
sine[2151] =494;
sine[2152] =494;
sine[2153] =494;
sine[2154] =495;
sine[2155] =495;
sine[2156] =495;
sine[2157] =495;
sine[2158] =495;
sine[2159] =495;
sine[2160] =495;
sine[2161] =496;
sine[2162] =496;
sine[2163] =496;
sine[2164] =496;
sine[2165] =496;
sine[2166] =496;
sine[2167] =496;
sine[2168] =496;
sine[2169] =497;
sine[2170] =497;
sine[2171] =497;
sine[2172] =497;
sine[2173] =497;
sine[2174] =497;
sine[2175] =497;
sine[2176] =497;
sine[2177] =498;
sine[2178] =498;
sine[2179] =498;
sine[2180] =498;
sine[2181] =498;
sine[2182] =498;
sine[2183] =498;
sine[2184] =498;
sine[2185] =499;
sine[2186] =499;
sine[2187] =499;
sine[2188] =499;
sine[2189] =499;
sine[2190] =499;
sine[2191] =499;
sine[2192] =499;
sine[2193] =500;
sine[2194] =500;
sine[2195] =500;
sine[2196] =500;
sine[2197] =500;
sine[2198] =500;
sine[2199] =500;
sine[2200] =500;
sine[2201] =500;
sine[2202] =501;
sine[2203] =501;
sine[2204] =501;
sine[2205] =501;
sine[2206] =501;
sine[2207] =501;
sine[2208] =501;
sine[2209] =501;
sine[2210] =501;
sine[2211] =502;
sine[2212] =502;
sine[2213] =502;
sine[2214] =502;
sine[2215] =502;
sine[2216] =502;
sine[2217] =502;
sine[2218] =502;
sine[2219] =502;
sine[2220] =502;
sine[2221] =503;
sine[2222] =503;
sine[2223] =503;
sine[2224] =503;
sine[2225] =503;
sine[2226] =503;
sine[2227] =503;
sine[2228] =503;
sine[2229] =503;
sine[2230] =503;
sine[2231] =504;
sine[2232] =504;
sine[2233] =504;
sine[2234] =504;
sine[2235] =504;
sine[2236] =504;
sine[2237] =504;
sine[2238] =504;
sine[2239] =504;
sine[2240] =504;
sine[2241] =504;
sine[2242] =505;
sine[2243] =505;
sine[2244] =505;
sine[2245] =505;
sine[2246] =505;
sine[2247] =505;
sine[2248] =505;
sine[2249] =505;
sine[2250] =505;
sine[2251] =505;
sine[2252] =505;
sine[2253] =505;
sine[2254] =506;
sine[2255] =506;
sine[2256] =506;
sine[2257] =506;
sine[2258] =506;
sine[2259] =506;
sine[2260] =506;
sine[2261] =506;
sine[2262] =506;
sine[2263] =506;
sine[2264] =506;
sine[2265] =506;
sine[2266] =506;
sine[2267] =507;
sine[2268] =507;
sine[2269] =507;
sine[2270] =507;
sine[2271] =507;
sine[2272] =507;
sine[2273] =507;
sine[2274] =507;
sine[2275] =507;
sine[2276] =507;
sine[2277] =507;
sine[2278] =507;
sine[2279] =507;
sine[2280] =507;
sine[2281] =508;
sine[2282] =508;
sine[2283] =508;
sine[2284] =508;
sine[2285] =508;
sine[2286] =508;
sine[2287] =508;
sine[2288] =508;
sine[2289] =508;
sine[2290] =508;
sine[2291] =508;
sine[2292] =508;
sine[2293] =508;
sine[2294] =508;
sine[2295] =508;
sine[2296] =508;
sine[2297] =508;
sine[2298] =509;
sine[2299] =509;
sine[2300] =509;
sine[2301] =509;
sine[2302] =509;
sine[2303] =509;
sine[2304] =509;
sine[2305] =509;
sine[2306] =509;
sine[2307] =509;
sine[2308] =509;
sine[2309] =509;
sine[2310] =509;
sine[2311] =509;
sine[2312] =509;
sine[2313] =509;
sine[2314] =509;
sine[2315] =509;
sine[2316] =509;
sine[2317] =509;
sine[2318] =509;
sine[2319] =510;
sine[2320] =510;
sine[2321] =510;
sine[2322] =510;
sine[2323] =510;
sine[2324] =510;
sine[2325] =510;
sine[2326] =510;
sine[2327] =510;
sine[2328] =510;
sine[2329] =510;
sine[2330] =510;
sine[2331] =510;
sine[2332] =510;
sine[2333] =510;
sine[2334] =510;
sine[2335] =510;
sine[2336] =510;
sine[2337] =510;
sine[2338] =510;
sine[2339] =510;
sine[2340] =510;
sine[2341] =510;
sine[2342] =510;
sine[2343] =510;
sine[2344] =510;
sine[2345] =510;
sine[2346] =510;
sine[2347] =510;
sine[2348] =510;
sine[2349] =511;
sine[2350] =511;
sine[2351] =511;
sine[2352] =511;
sine[2353] =511;
sine[2354] =511;
sine[2355] =511;
sine[2356] =511;
sine[2357] =511;
sine[2358] =511;
sine[2359] =511;
sine[2360] =511;
sine[2361] =511;
sine[2362] =511;
sine[2363] =511;
sine[2364] =511;
sine[2365] =511;
sine[2366] =511;
sine[2367] =511;
sine[2368] =511;
sine[2369] =511;
sine[2370] =511;
sine[2371] =511;
sine[2372] =511;
sine[2373] =511;
sine[2374] =511;
sine[2375] =511;
sine[2376] =511;
sine[2377] =511;
sine[2378] =511;
sine[2379] =511;
sine[2380] =511;
sine[2381] =511;
sine[2382] =511;
sine[2383] =511;
sine[2384] =511;
sine[2385] =511;
sine[2386] =511;
sine[2387] =511;
sine[2388] =511;
sine[2389] =511;
sine[2390] =511;
sine[2391] =511;
sine[2392] =511;
sine[2393] =511;
sine[2394] =511;
sine[2395] =511;
sine[2396] =511;
sine[2397] =511;
sine[2398] =511;
sine[2399] =511;
sine[2400] =511;
sine[2401] =511;
sine[2402] =511;
sine[2403] =511;
sine[2404] =511;
sine[2405] =511;
sine[2406] =511;
sine[2407] =511;
sine[2408] =511;
sine[2409] =511;
sine[2410] =511;
sine[2411] =511;
sine[2412] =511;
sine[2413] =511;
sine[2414] =511;
sine[2415] =511;
sine[2416] =511;
sine[2417] =511;
sine[2418] =511;
sine[2419] =511;
sine[2420] =511;
sine[2421] =511;
sine[2422] =511;
sine[2423] =511;
sine[2424] =511;
sine[2425] =511;
sine[2426] =511;
sine[2427] =511;
sine[2428] =511;
sine[2429] =511;
sine[2430] =510;
sine[2431] =510;
sine[2432] =510;
sine[2433] =510;
sine[2434] =510;
sine[2435] =510;
sine[2436] =510;
sine[2437] =510;
sine[2438] =510;
sine[2439] =510;
sine[2440] =510;
sine[2441] =510;
sine[2442] =510;
sine[2443] =510;
sine[2444] =510;
sine[2445] =510;
sine[2446] =510;
sine[2447] =510;
sine[2448] =510;
sine[2449] =510;
sine[2450] =510;
sine[2451] =510;
sine[2452] =510;
sine[2453] =510;
sine[2454] =510;
sine[2455] =510;
sine[2456] =510;
sine[2457] =510;
sine[2458] =510;
sine[2459] =510;
sine[2460] =509;
sine[2461] =509;
sine[2462] =509;
sine[2463] =509;
sine[2464] =509;
sine[2465] =509;
sine[2466] =509;
sine[2467] =509;
sine[2468] =509;
sine[2469] =509;
sine[2470] =509;
sine[2471] =509;
sine[2472] =509;
sine[2473] =509;
sine[2474] =509;
sine[2475] =509;
sine[2476] =509;
sine[2477] =509;
sine[2478] =509;
sine[2479] =509;
sine[2480] =509;
sine[2481] =508;
sine[2482] =508;
sine[2483] =508;
sine[2484] =508;
sine[2485] =508;
sine[2486] =508;
sine[2487] =508;
sine[2488] =508;
sine[2489] =508;
sine[2490] =508;
sine[2491] =508;
sine[2492] =508;
sine[2493] =508;
sine[2494] =508;
sine[2495] =508;
sine[2496] =508;
sine[2497] =508;
sine[2498] =507;
sine[2499] =507;
sine[2500] =507;
sine[2501] =507;
sine[2502] =507;
sine[2503] =507;
sine[2504] =507;
sine[2505] =507;
sine[2506] =507;
sine[2507] =507;
sine[2508] =507;
sine[2509] =507;
sine[2510] =507;
sine[2511] =507;
sine[2512] =506;
sine[2513] =506;
sine[2514] =506;
sine[2515] =506;
sine[2516] =506;
sine[2517] =506;
sine[2518] =506;
sine[2519] =506;
sine[2520] =506;
sine[2521] =506;
sine[2522] =506;
sine[2523] =506;
sine[2524] =506;
sine[2525] =505;
sine[2526] =505;
sine[2527] =505;
sine[2528] =505;
sine[2529] =505;
sine[2530] =505;
sine[2531] =505;
sine[2532] =505;
sine[2533] =505;
sine[2534] =505;
sine[2535] =505;
sine[2536] =505;
sine[2537] =504;
sine[2538] =504;
sine[2539] =504;
sine[2540] =504;
sine[2541] =504;
sine[2542] =504;
sine[2543] =504;
sine[2544] =504;
sine[2545] =504;
sine[2546] =504;
sine[2547] =504;
sine[2548] =503;
sine[2549] =503;
sine[2550] =503;
sine[2551] =503;
sine[2552] =503;
sine[2553] =503;
sine[2554] =503;
sine[2555] =503;
sine[2556] =503;
sine[2557] =503;
sine[2558] =502;
sine[2559] =502;
sine[2560] =502;
sine[2561] =502;
sine[2562] =502;
sine[2563] =502;
sine[2564] =502;
sine[2565] =502;
sine[2566] =502;
sine[2567] =502;
sine[2568] =501;
sine[2569] =501;
sine[2570] =501;
sine[2571] =501;
sine[2572] =501;
sine[2573] =501;
sine[2574] =501;
sine[2575] =501;
sine[2576] =501;
sine[2577] =500;
sine[2578] =500;
sine[2579] =500;
sine[2580] =500;
sine[2581] =500;
sine[2582] =500;
sine[2583] =500;
sine[2584] =500;
sine[2585] =500;
sine[2586] =499;
sine[2587] =499;
sine[2588] =499;
sine[2589] =499;
sine[2590] =499;
sine[2591] =499;
sine[2592] =499;
sine[2593] =499;
sine[2594] =498;
sine[2595] =498;
sine[2596] =498;
sine[2597] =498;
sine[2598] =498;
sine[2599] =498;
sine[2600] =498;
sine[2601] =498;
sine[2602] =497;
sine[2603] =497;
sine[2604] =497;
sine[2605] =497;
sine[2606] =497;
sine[2607] =497;
sine[2608] =497;
sine[2609] =497;
sine[2610] =496;
sine[2611] =496;
sine[2612] =496;
sine[2613] =496;
sine[2614] =496;
sine[2615] =496;
sine[2616] =496;
sine[2617] =496;
sine[2618] =495;
sine[2619] =495;
sine[2620] =495;
sine[2621] =495;
sine[2622] =495;
sine[2623] =495;
sine[2624] =495;
sine[2625] =494;
sine[2626] =494;
sine[2627] =494;
sine[2628] =494;
sine[2629] =494;
sine[2630] =494;
sine[2631] =494;
sine[2632] =493;
sine[2633] =493;
sine[2634] =493;
sine[2635] =493;
sine[2636] =493;
sine[2637] =493;
sine[2638] =493;
sine[2639] =492;
sine[2640] =492;
sine[2641] =492;
sine[2642] =492;
sine[2643] =492;
sine[2644] =492;
sine[2645] =492;
sine[2646] =491;
sine[2647] =491;
sine[2648] =491;
sine[2649] =491;
sine[2650] =491;
sine[2651] =491;
sine[2652] =490;
sine[2653] =490;
sine[2654] =490;
sine[2655] =490;
sine[2656] =490;
sine[2657] =490;
sine[2658] =490;
sine[2659] =489;
sine[2660] =489;
sine[2661] =489;
sine[2662] =489;
sine[2663] =489;
sine[2664] =489;
sine[2665] =488;
sine[2666] =488;
sine[2667] =488;
sine[2668] =488;
sine[2669] =488;
sine[2670] =488;
sine[2671] =487;
sine[2672] =487;
sine[2673] =487;
sine[2674] =487;
sine[2675] =487;
sine[2676] =487;
sine[2677] =486;
sine[2678] =486;
sine[2679] =486;
sine[2680] =486;
sine[2681] =486;
sine[2682] =486;
sine[2683] =485;
sine[2684] =485;
sine[2685] =485;
sine[2686] =485;
sine[2687] =485;
sine[2688] =485;
sine[2689] =484;
sine[2690] =484;
sine[2691] =484;
sine[2692] =484;
sine[2693] =484;
sine[2694] =484;
sine[2695] =483;
sine[2696] =483;
sine[2697] =483;
sine[2698] =483;
sine[2699] =483;
sine[2700] =482;
sine[2701] =482;
sine[2702] =482;
sine[2703] =482;
sine[2704] =482;
sine[2705] =482;
sine[2706] =481;
sine[2707] =481;
sine[2708] =481;
sine[2709] =481;
sine[2710] =481;
sine[2711] =480;
sine[2712] =480;
sine[2713] =480;
sine[2714] =480;
sine[2715] =480;
sine[2716] =480;
sine[2717] =479;
sine[2718] =479;
sine[2719] =479;
sine[2720] =479;
sine[2721] =479;
sine[2722] =478;
sine[2723] =478;
sine[2724] =478;
sine[2725] =478;
sine[2726] =478;
sine[2727] =477;
sine[2728] =477;
sine[2729] =477;
sine[2730] =477;
sine[2731] =477;
sine[2732] =476;
sine[2733] =476;
sine[2734] =476;
sine[2735] =476;
sine[2736] =476;
sine[2737] =475;
sine[2738] =475;
sine[2739] =475;
sine[2740] =475;
sine[2741] =475;
sine[2742] =474;
sine[2743] =474;
sine[2744] =474;
sine[2745] =474;
sine[2746] =474;
sine[2747] =473;
sine[2748] =473;
sine[2749] =473;
sine[2750] =473;
sine[2751] =473;
sine[2752] =472;
sine[2753] =472;
sine[2754] =472;
sine[2755] =472;
sine[2756] =472;
sine[2757] =471;
sine[2758] =471;
sine[2759] =471;
sine[2760] =471;
sine[2761] =471;
sine[2762] =470;
sine[2763] =470;
sine[2764] =470;
sine[2765] =470;
sine[2766] =469;
sine[2767] =469;
sine[2768] =469;
sine[2769] =469;
sine[2770] =469;
sine[2771] =468;
sine[2772] =468;
sine[2773] =468;
sine[2774] =468;
sine[2775] =468;
sine[2776] =467;
sine[2777] =467;
sine[2778] =467;
sine[2779] =467;
sine[2780] =466;
sine[2781] =466;
sine[2782] =466;
sine[2783] =466;
sine[2784] =466;
sine[2785] =465;
sine[2786] =465;
sine[2787] =465;
sine[2788] =465;
sine[2789] =464;
sine[2790] =464;
sine[2791] =464;
sine[2792] =464;
sine[2793] =463;
sine[2794] =463;
sine[2795] =463;
sine[2796] =463;
sine[2797] =463;
sine[2798] =462;
sine[2799] =462;
sine[2800] =462;
sine[2801] =462;
sine[2802] =461;
sine[2803] =461;
sine[2804] =461;
sine[2805] =461;
sine[2806] =460;
sine[2807] =460;
sine[2808] =460;
sine[2809] =460;
sine[2810] =460;
sine[2811] =459;
sine[2812] =459;
sine[2813] =459;
sine[2814] =459;
sine[2815] =458;
sine[2816] =458;
sine[2817] =458;
sine[2818] =458;
sine[2819] =457;
sine[2820] =457;
sine[2821] =457;
sine[2822] =457;
sine[2823] =456;
sine[2824] =456;
sine[2825] =456;
sine[2826] =456;
sine[2827] =455;
sine[2828] =455;
sine[2829] =455;
sine[2830] =455;
sine[2831] =454;
sine[2832] =454;
sine[2833] =454;
sine[2834] =454;
sine[2835] =454;
sine[2836] =453;
sine[2837] =453;
sine[2838] =453;
sine[2839] =453;
sine[2840] =452;
sine[2841] =452;
sine[2842] =452;
sine[2843] =452;
sine[2844] =451;
sine[2845] =451;
sine[2846] =451;
sine[2847] =450;
sine[2848] =450;
sine[2849] =450;
sine[2850] =450;
sine[2851] =449;
sine[2852] =449;
sine[2853] =449;
sine[2854] =449;
sine[2855] =448;
sine[2856] =448;
sine[2857] =448;
sine[2858] =448;
sine[2859] =447;
sine[2860] =447;
sine[2861] =447;
sine[2862] =447;
sine[2863] =446;
sine[2864] =446;
sine[2865] =446;
sine[2866] =446;
sine[2867] =445;
sine[2868] =445;
sine[2869] =445;
sine[2870] =445;
sine[2871] =444;
sine[2872] =444;
sine[2873] =444;
sine[2874] =443;
sine[2875] =443;
sine[2876] =443;
sine[2877] =443;
sine[2878] =442;
sine[2879] =442;
sine[2880] =442;
sine[2881] =442;
sine[2882] =441;
sine[2883] =441;
sine[2884] =441;
sine[2885] =441;
sine[2886] =440;
sine[2887] =440;
sine[2888] =440;
sine[2889] =439;
sine[2890] =439;
sine[2891] =439;
sine[2892] =439;
sine[2893] =438;
sine[2894] =438;
sine[2895] =438;
sine[2896] =438;
sine[2897] =437;
sine[2898] =437;
sine[2899] =437;
sine[2900] =436;
sine[2901] =436;
sine[2902] =436;
sine[2903] =436;
sine[2904] =435;
sine[2905] =435;
sine[2906] =435;
sine[2907] =434;
sine[2908] =434;
sine[2909] =434;
sine[2910] =434;
sine[2911] =433;
sine[2912] =433;
sine[2913] =433;
sine[2914] =433;
sine[2915] =432;
sine[2916] =432;
sine[2917] =432;
sine[2918] =431;
sine[2919] =431;
sine[2920] =431;
sine[2921] =431;
sine[2922] =430;
sine[2923] =430;
sine[2924] =430;
sine[2925] =429;
sine[2926] =429;
sine[2927] =429;
sine[2928] =429;
sine[2929] =428;
sine[2930] =428;
sine[2931] =428;
sine[2932] =427;
sine[2933] =427;
sine[2934] =427;
sine[2935] =427;
sine[2936] =426;
sine[2937] =426;
sine[2938] =426;
sine[2939] =425;
sine[2940] =425;
sine[2941] =425;
sine[2942] =424;
sine[2943] =424;
sine[2944] =424;
sine[2945] =424;
sine[2946] =423;
sine[2947] =423;
sine[2948] =423;
sine[2949] =422;
sine[2950] =422;
sine[2951] =422;
sine[2952] =421;
sine[2953] =421;
sine[2954] =421;
sine[2955] =421;
sine[2956] =420;
sine[2957] =420;
sine[2958] =420;
sine[2959] =419;
sine[2960] =419;
sine[2961] =419;
sine[2962] =418;
sine[2963] =418;
sine[2964] =418;
sine[2965] =418;
sine[2966] =417;
sine[2967] =417;
sine[2968] =417;
sine[2969] =416;
sine[2970] =416;
sine[2971] =416;
sine[2972] =415;
sine[2973] =415;
sine[2974] =415;
sine[2975] =415;
sine[2976] =414;
sine[2977] =414;
sine[2978] =414;
sine[2979] =413;
sine[2980] =413;
sine[2981] =413;
sine[2982] =412;
sine[2983] =412;
sine[2984] =412;
sine[2985] =411;
sine[2986] =411;
sine[2987] =411;
sine[2988] =411;
sine[2989] =410;
sine[2990] =410;
sine[2991] =410;
sine[2992] =409;
sine[2993] =409;
sine[2994] =409;
sine[2995] =408;
sine[2996] =408;
sine[2997] =408;
sine[2998] =407;
sine[2999] =407;
sine[3000] =407;
sine[3001] =406;
sine[3002] =406;
sine[3003] =406;
sine[3004] =405;
sine[3005] =405;
sine[3006] =405;
sine[3007] =405;
sine[3008] =404;
sine[3009] =404;
sine[3010] =404;
sine[3011] =403;
sine[3012] =403;
sine[3013] =403;
sine[3014] =402;
sine[3015] =402;
sine[3016] =402;
sine[3017] =401;
sine[3018] =401;
sine[3019] =401;
sine[3020] =400;
sine[3021] =400;
sine[3022] =400;
sine[3023] =399;
sine[3024] =399;
sine[3025] =399;
sine[3026] =398;
sine[3027] =398;
sine[3028] =398;
sine[3029] =397;
sine[3030] =397;
sine[3031] =397;
sine[3032] =396;
sine[3033] =396;
sine[3034] =396;
sine[3035] =395;
sine[3036] =395;
sine[3037] =395;
sine[3038] =395;
sine[3039] =394;
sine[3040] =394;
sine[3041] =394;
sine[3042] =393;
sine[3043] =393;
sine[3044] =393;
sine[3045] =392;
sine[3046] =392;
sine[3047] =392;
sine[3048] =391;
sine[3049] =391;
sine[3050] =391;
sine[3051] =390;
sine[3052] =390;
sine[3053] =390;
sine[3054] =389;
sine[3055] =389;
sine[3056] =389;
sine[3057] =388;
sine[3058] =388;
sine[3059] =388;
sine[3060] =387;
sine[3061] =387;
sine[3062] =387;
sine[3063] =386;
sine[3064] =386;
sine[3065] =386;
sine[3066] =385;
sine[3067] =385;
sine[3068] =384;
sine[3069] =384;
sine[3070] =384;
sine[3071] =383;
sine[3072] =383;
sine[3073] =383;
sine[3074] =382;
sine[3075] =382;
sine[3076] =382;
sine[3077] =381;
sine[3078] =381;
sine[3079] =381;
sine[3080] =380;
sine[3081] =380;
sine[3082] =380;
sine[3083] =379;
sine[3084] =379;
sine[3085] =379;
sine[3086] =378;
sine[3087] =378;
sine[3088] =378;
sine[3089] =377;
sine[3090] =377;
sine[3091] =377;
sine[3092] =376;
sine[3093] =376;
sine[3094] =376;
sine[3095] =375;
sine[3096] =375;
sine[3097] =375;
sine[3098] =374;
sine[3099] =374;
sine[3100] =374;
sine[3101] =373;
sine[3102] =373;
sine[3103] =372;
sine[3104] =372;
sine[3105] =372;
sine[3106] =371;
sine[3107] =371;
sine[3108] =371;
sine[3109] =370;
sine[3110] =370;
sine[3111] =370;
sine[3112] =369;
sine[3113] =369;
sine[3114] =369;
sine[3115] =368;
sine[3116] =368;
sine[3117] =368;
sine[3118] =367;
sine[3119] =367;
sine[3120] =367;
sine[3121] =366;
sine[3122] =366;
sine[3123] =365;
sine[3124] =365;
sine[3125] =365;
sine[3126] =364;
sine[3127] =364;
sine[3128] =364;
sine[3129] =363;
sine[3130] =363;
sine[3131] =363;
sine[3132] =362;
sine[3133] =362;
sine[3134] =362;
sine[3135] =361;
sine[3136] =361;
sine[3137] =360;
sine[3138] =360;
sine[3139] =360;
sine[3140] =359;
sine[3141] =359;
sine[3142] =359;
sine[3143] =358;
sine[3144] =358;
sine[3145] =358;
sine[3146] =357;
sine[3147] =357;
sine[3148] =357;
sine[3149] =356;
sine[3150] =356;
sine[3151] =355;
sine[3152] =355;
sine[3153] =355;
sine[3154] =354;
sine[3155] =354;
sine[3156] =354;
sine[3157] =353;
sine[3158] =353;
sine[3159] =353;
sine[3160] =352;
sine[3161] =352;
sine[3162] =351;
sine[3163] =351;
sine[3164] =351;
sine[3165] =350;
sine[3166] =350;
sine[3167] =350;
sine[3168] =349;
sine[3169] =349;
sine[3170] =349;
sine[3171] =348;
sine[3172] =348;
sine[3173] =347;
sine[3174] =347;
sine[3175] =347;
sine[3176] =346;
sine[3177] =346;
sine[3178] =346;
sine[3179] =345;
sine[3180] =345;
sine[3181] =345;
sine[3182] =344;
sine[3183] =344;
sine[3184] =343;
sine[3185] =343;
sine[3186] =343;
sine[3187] =342;
sine[3188] =342;
sine[3189] =342;
sine[3190] =341;
sine[3191] =341;
sine[3192] =340;
sine[3193] =340;
sine[3194] =340;
sine[3195] =339;
sine[3196] =339;
sine[3197] =339;
sine[3198] =338;
sine[3199] =338;
sine[3200] =338;
sine[3201] =337;
sine[3202] =337;
sine[3203] =336;
sine[3204] =336;
sine[3205] =336;
sine[3206] =335;
sine[3207] =335;
sine[3208] =335;
sine[3209] =334;
sine[3210] =334;
sine[3211] =333;
sine[3212] =333;
sine[3213] =333;
sine[3214] =332;
sine[3215] =332;
sine[3216] =332;
sine[3217] =331;
sine[3218] =331;
sine[3219] =330;
sine[3220] =330;
sine[3221] =330;
sine[3222] =329;
sine[3223] =329;
sine[3224] =329;
sine[3225] =328;
sine[3226] =328;
sine[3227] =327;
sine[3228] =327;
sine[3229] =327;
sine[3230] =326;
sine[3231] =326;
sine[3232] =326;
sine[3233] =325;
sine[3234] =325;
sine[3235] =324;
sine[3236] =324;
sine[3237] =324;
sine[3238] =323;
sine[3239] =323;
sine[3240] =323;
sine[3241] =322;
sine[3242] =322;
sine[3243] =321;
sine[3244] =321;
sine[3245] =321;
sine[3246] =320;
sine[3247] =320;
sine[3248] =319;
sine[3249] =319;
sine[3250] =319;
sine[3251] =318;
sine[3252] =318;
sine[3253] =318;
sine[3254] =317;
sine[3255] =317;
sine[3256] =316;
sine[3257] =316;
sine[3258] =316;
sine[3259] =315;
sine[3260] =315;
sine[3261] =315;
sine[3262] =314;
sine[3263] =314;
sine[3264] =313;
sine[3265] =313;
sine[3266] =313;
sine[3267] =312;
sine[3268] =312;
sine[3269] =311;
sine[3270] =311;
sine[3271] =311;
sine[3272] =310;
sine[3273] =310;
sine[3274] =310;
sine[3275] =309;
sine[3276] =309;
sine[3277] =308;
sine[3278] =308;
sine[3279] =308;
sine[3280] =307;
sine[3281] =307;
sine[3282] =306;
sine[3283] =306;
sine[3284] =306;
sine[3285] =305;
sine[3286] =305;
sine[3287] =305;
sine[3288] =304;
sine[3289] =304;
sine[3290] =303;
sine[3291] =303;
sine[3292] =303;
sine[3293] =302;
sine[3294] =302;
sine[3295] =301;
sine[3296] =301;
sine[3297] =301;
sine[3298] =300;
sine[3299] =300;
sine[3300] =300;
sine[3301] =299;
sine[3302] =299;
sine[3303] =298;
sine[3304] =298;
sine[3305] =298;
sine[3306] =297;
sine[3307] =297;
sine[3308] =296;
sine[3309] =296;
sine[3310] =296;
sine[3311] =295;
sine[3312] =295;
sine[3313] =295;
sine[3314] =294;
sine[3315] =294;
sine[3316] =293;
sine[3317] =293;
sine[3318] =293;
sine[3319] =292;
sine[3320] =292;
sine[3321] =291;
sine[3322] =291;
sine[3323] =291;
sine[3324] =290;
sine[3325] =290;
sine[3326] =289;
sine[3327] =289;
sine[3328] =289;
sine[3329] =288;
sine[3330] =288;
sine[3331] =288;
sine[3332] =287;
sine[3333] =287;
sine[3334] =286;
sine[3335] =286;
sine[3336] =286;
sine[3337] =285;
sine[3338] =285;
sine[3339] =284;
sine[3340] =284;
sine[3341] =284;
sine[3342] =283;
sine[3343] =283;
sine[3344] =282;
sine[3345] =282;
sine[3346] =282;
sine[3347] =281;
sine[3348] =281;
sine[3349] =281;
sine[3350] =280;
sine[3351] =280;
sine[3352] =279;
sine[3353] =279;
sine[3354] =279;
sine[3355] =278;
sine[3356] =278;
sine[3357] =277;
sine[3358] =277;
sine[3359] =277;
sine[3360] =276;
sine[3361] =276;
sine[3362] =275;
sine[3363] =275;
sine[3364] =275;
sine[3365] =274;
sine[3366] =274;
sine[3367] =274;
sine[3368] =273;
sine[3369] =273;
sine[3370] =272;
sine[3371] =272;
sine[3372] =272;
sine[3373] =271;
sine[3374] =271;
sine[3375] =270;
sine[3376] =270;
sine[3377] =270;
sine[3378] =269;
sine[3379] =269;
sine[3380] =268;
sine[3381] =268;
sine[3382] =268;
sine[3383] =267;
sine[3384] =267;
sine[3385] =266;
sine[3386] =266;
sine[3387] =266;
sine[3388] =265;
sine[3389] =265;
sine[3390] =265;
sine[3391] =264;
sine[3392] =264;
sine[3393] =263;
sine[3394] =263;
sine[3395] =263;
sine[3396] =262;
sine[3397] =262;
sine[3398] =261;
sine[3399] =261;
sine[3400] =261;
sine[3401] =260;
sine[3402] =260;
sine[3403] =259;
sine[3404] =259;
sine[3405] =259;
sine[3406] =258;
sine[3407] =258;
sine[3408] =257;
sine[3409] =257;
sine[3410] =257;
sine[3411] =256;
sine[3412] =256;
sine[3413] =256;
sine[3414] =255;
sine[3415] =255;
sine[3416] =254;
sine[3417] =254;
sine[3418] =254;
sine[3419] =253;
sine[3420] =253;
sine[3421] =252;
sine[3422] =252;
sine[3423] =252;
sine[3424] =251;
sine[3425] =251;
sine[3426] =250;
sine[3427] =250;
sine[3428] =250;
sine[3429] =249;
sine[3430] =249;
sine[3431] =248;
sine[3432] =248;
sine[3433] =248;
sine[3434] =247;
sine[3435] =247;
sine[3436] =246;
sine[3437] =246;
sine[3438] =246;
sine[3439] =245;
sine[3440] =245;
sine[3441] =245;
sine[3442] =244;
sine[3443] =244;
sine[3444] =243;
sine[3445] =243;
sine[3446] =243;
sine[3447] =242;
sine[3448] =242;
sine[3449] =241;
sine[3450] =241;
sine[3451] =241;
sine[3452] =240;
sine[3453] =240;
sine[3454] =239;
sine[3455] =239;
sine[3456] =239;
sine[3457] =238;
sine[3458] =238;
sine[3459] =237;
sine[3460] =237;
sine[3461] =237;
sine[3462] =236;
sine[3463] =236;
sine[3464] =236;
sine[3465] =235;
sine[3466] =235;
sine[3467] =234;
sine[3468] =234;
sine[3469] =234;
sine[3470] =233;
sine[3471] =233;
sine[3472] =232;
sine[3473] =232;
sine[3474] =232;
sine[3475] =231;
sine[3476] =231;
sine[3477] =230;
sine[3478] =230;
sine[3479] =230;
sine[3480] =229;
sine[3481] =229;
sine[3482] =229;
sine[3483] =228;
sine[3484] =228;
sine[3485] =227;
sine[3486] =227;
sine[3487] =227;
sine[3488] =226;
sine[3489] =226;
sine[3490] =225;
sine[3491] =225;
sine[3492] =225;
sine[3493] =224;
sine[3494] =224;
sine[3495] =223;
sine[3496] =223;
sine[3497] =223;
sine[3498] =222;
sine[3499] =222;
sine[3500] =222;
sine[3501] =221;
sine[3502] =221;
sine[3503] =220;
sine[3504] =220;
sine[3505] =220;
sine[3506] =219;
sine[3507] =219;
sine[3508] =218;
sine[3509] =218;
sine[3510] =218;
sine[3511] =217;
sine[3512] =217;
sine[3513] =216;
sine[3514] =216;
sine[3515] =216;
sine[3516] =215;
sine[3517] =215;
sine[3518] =215;
sine[3519] =214;
sine[3520] =214;
sine[3521] =213;
sine[3522] =213;
sine[3523] =213;
sine[3524] =212;
sine[3525] =212;
sine[3526] =211;
sine[3527] =211;
sine[3528] =211;
sine[3529] =210;
sine[3530] =210;
sine[3531] =210;
sine[3532] =209;
sine[3533] =209;
sine[3534] =208;
sine[3535] =208;
sine[3536] =208;
sine[3537] =207;
sine[3538] =207;
sine[3539] =206;
sine[3540] =206;
sine[3541] =206;
sine[3542] =205;
sine[3543] =205;
sine[3544] =205;
sine[3545] =204;
sine[3546] =204;
sine[3547] =203;
sine[3548] =203;
sine[3549] =203;
sine[3550] =202;
sine[3551] =202;
sine[3552] =201;
sine[3553] =201;
sine[3554] =201;
sine[3555] =200;
sine[3556] =200;
sine[3557] =200;
sine[3558] =199;
sine[3559] =199;
sine[3560] =198;
sine[3561] =198;
sine[3562] =198;
sine[3563] =197;
sine[3564] =197;
sine[3565] =196;
sine[3566] =196;
sine[3567] =196;
sine[3568] =195;
sine[3569] =195;
sine[3570] =195;
sine[3571] =194;
sine[3572] =194;
sine[3573] =193;
sine[3574] =193;
sine[3575] =193;
sine[3576] =192;
sine[3577] =192;
sine[3578] =192;
sine[3579] =191;
sine[3580] =191;
sine[3581] =190;
sine[3582] =190;
sine[3583] =190;
sine[3584] =189;
sine[3585] =189;
sine[3586] =188;
sine[3587] =188;
sine[3588] =188;
sine[3589] =187;
sine[3590] =187;
sine[3591] =187;
sine[3592] =186;
sine[3593] =186;
sine[3594] =185;
sine[3595] =185;
sine[3596] =185;
sine[3597] =184;
sine[3598] =184;
sine[3599] =184;
sine[3600] =183;
sine[3601] =183;
sine[3602] =182;
sine[3603] =182;
sine[3604] =182;
sine[3605] =181;
sine[3606] =181;
sine[3607] =181;
sine[3608] =180;
sine[3609] =180;
sine[3610] =179;
sine[3611] =179;
sine[3612] =179;
sine[3613] =178;
sine[3614] =178;
sine[3615] =178;
sine[3616] =177;
sine[3617] =177;
sine[3618] =176;
sine[3619] =176;
sine[3620] =176;
sine[3621] =175;
sine[3622] =175;
sine[3623] =175;
sine[3624] =174;
sine[3625] =174;
sine[3626] =173;
sine[3627] =173;
sine[3628] =173;
sine[3629] =172;
sine[3630] =172;
sine[3631] =172;
sine[3632] =171;
sine[3633] =171;
sine[3634] =171;
sine[3635] =170;
sine[3636] =170;
sine[3637] =169;
sine[3638] =169;
sine[3639] =169;
sine[3640] =168;
sine[3641] =168;
sine[3642] =168;
sine[3643] =167;
sine[3644] =167;
sine[3645] =166;
sine[3646] =166;
sine[3647] =166;
sine[3648] =165;
sine[3649] =165;
sine[3650] =165;
sine[3651] =164;
sine[3652] =164;
sine[3653] =164;
sine[3654] =163;
sine[3655] =163;
sine[3656] =162;
sine[3657] =162;
sine[3658] =162;
sine[3659] =161;
sine[3660] =161;
sine[3661] =161;
sine[3662] =160;
sine[3663] =160;
sine[3664] =160;
sine[3665] =159;
sine[3666] =159;
sine[3667] =158;
sine[3668] =158;
sine[3669] =158;
sine[3670] =157;
sine[3671] =157;
sine[3672] =157;
sine[3673] =156;
sine[3674] =156;
sine[3675] =156;
sine[3676] =155;
sine[3677] =155;
sine[3678] =154;
sine[3679] =154;
sine[3680] =154;
sine[3681] =153;
sine[3682] =153;
sine[3683] =153;
sine[3684] =152;
sine[3685] =152;
sine[3686] =152;
sine[3687] =151;
sine[3688] =151;
sine[3689] =151;
sine[3690] =150;
sine[3691] =150;
sine[3692] =149;
sine[3693] =149;
sine[3694] =149;
sine[3695] =148;
sine[3696] =148;
sine[3697] =148;
sine[3698] =147;
sine[3699] =147;
sine[3700] =147;
sine[3701] =146;
sine[3702] =146;
sine[3703] =146;
sine[3704] =145;
sine[3705] =145;
sine[3706] =144;
sine[3707] =144;
sine[3708] =144;
sine[3709] =143;
sine[3710] =143;
sine[3711] =143;
sine[3712] =142;
sine[3713] =142;
sine[3714] =142;
sine[3715] =141;
sine[3716] =141;
sine[3717] =141;
sine[3718] =140;
sine[3719] =140;
sine[3720] =140;
sine[3721] =139;
sine[3722] =139;
sine[3723] =139;
sine[3724] =138;
sine[3725] =138;
sine[3726] =137;
sine[3727] =137;
sine[3728] =137;
sine[3729] =136;
sine[3730] =136;
sine[3731] =136;
sine[3732] =135;
sine[3733] =135;
sine[3734] =135;
sine[3735] =134;
sine[3736] =134;
sine[3737] =134;
sine[3738] =133;
sine[3739] =133;
sine[3740] =133;
sine[3741] =132;
sine[3742] =132;
sine[3743] =132;
sine[3744] =131;
sine[3745] =131;
sine[3746] =131;
sine[3747] =130;
sine[3748] =130;
sine[3749] =130;
sine[3750] =129;
sine[3751] =129;
sine[3752] =129;
sine[3753] =128;
sine[3754] =128;
sine[3755] =128;
sine[3756] =127;
sine[3757] =127;
sine[3758] =127;
sine[3759] =126;
sine[3760] =126;
sine[3761] =125;
sine[3762] =125;
sine[3763] =125;
sine[3764] =124;
sine[3765] =124;
sine[3766] =124;
sine[3767] =123;
sine[3768] =123;
sine[3769] =123;
sine[3770] =122;
sine[3771] =122;
sine[3772] =122;
sine[3773] =121;
sine[3774] =121;
sine[3775] =121;
sine[3776] =120;
sine[3777] =120;
sine[3778] =120;
sine[3779] =119;
sine[3780] =119;
sine[3781] =119;
sine[3782] =118;
sine[3783] =118;
sine[3784] =118;
sine[3785] =117;
sine[3786] =117;
sine[3787] =117;
sine[3788] =116;
sine[3789] =116;
sine[3790] =116;
sine[3791] =116;
sine[3792] =115;
sine[3793] =115;
sine[3794] =115;
sine[3795] =114;
sine[3796] =114;
sine[3797] =114;
sine[3798] =113;
sine[3799] =113;
sine[3800] =113;
sine[3801] =112;
sine[3802] =112;
sine[3803] =112;
sine[3804] =111;
sine[3805] =111;
sine[3806] =111;
sine[3807] =110;
sine[3808] =110;
sine[3809] =110;
sine[3810] =109;
sine[3811] =109;
sine[3812] =109;
sine[3813] =108;
sine[3814] =108;
sine[3815] =108;
sine[3816] =107;
sine[3817] =107;
sine[3818] =107;
sine[3819] =106;
sine[3820] =106;
sine[3821] =106;
sine[3822] =106;
sine[3823] =105;
sine[3824] =105;
sine[3825] =105;
sine[3826] =104;
sine[3827] =104;
sine[3828] =104;
sine[3829] =103;
sine[3830] =103;
sine[3831] =103;
sine[3832] =102;
sine[3833] =102;
sine[3834] =102;
sine[3835] =101;
sine[3836] =101;
sine[3837] =101;
sine[3838] =100;
sine[3839] =100;
sine[3840] =100;
sine[3841] =100;
sine[3842] =99;
sine[3843] =99;
sine[3844] =99;
sine[3845] =98;
sine[3846] =98;
sine[3847] =98;
sine[3848] =97;
sine[3849] =97;
sine[3850] =97;
sine[3851] =96;
sine[3852] =96;
sine[3853] =96;
sine[3854] =96;
sine[3855] =95;
sine[3856] =95;
sine[3857] =95;
sine[3858] =94;
sine[3859] =94;
sine[3860] =94;
sine[3861] =93;
sine[3862] =93;
sine[3863] =93;
sine[3864] =93;
sine[3865] =92;
sine[3866] =92;
sine[3867] =92;
sine[3868] =91;
sine[3869] =91;
sine[3870] =91;
sine[3871] =90;
sine[3872] =90;
sine[3873] =90;
sine[3874] =90;
sine[3875] =89;
sine[3876] =89;
sine[3877] =89;
sine[3878] =88;
sine[3879] =88;
sine[3880] =88;
sine[3881] =87;
sine[3882] =87;
sine[3883] =87;
sine[3884] =87;
sine[3885] =86;
sine[3886] =86;
sine[3887] =86;
sine[3888] =85;
sine[3889] =85;
sine[3890] =85;
sine[3891] =84;
sine[3892] =84;
sine[3893] =84;
sine[3894] =84;
sine[3895] =83;
sine[3896] =83;
sine[3897] =83;
sine[3898] =82;
sine[3899] =82;
sine[3900] =82;
sine[3901] =82;
sine[3902] =81;
sine[3903] =81;
sine[3904] =81;
sine[3905] =80;
sine[3906] =80;
sine[3907] =80;
sine[3908] =80;
sine[3909] =79;
sine[3910] =79;
sine[3911] =79;
sine[3912] =78;
sine[3913] =78;
sine[3914] =78;
sine[3915] =78;
sine[3916] =77;
sine[3917] =77;
sine[3918] =77;
sine[3919] =77;
sine[3920] =76;
sine[3921] =76;
sine[3922] =76;
sine[3923] =75;
sine[3924] =75;
sine[3925] =75;
sine[3926] =75;
sine[3927] =74;
sine[3928] =74;
sine[3929] =74;
sine[3930] =73;
sine[3931] =73;
sine[3932] =73;
sine[3933] =73;
sine[3934] =72;
sine[3935] =72;
sine[3936] =72;
sine[3937] =72;
sine[3938] =71;
sine[3939] =71;
sine[3940] =71;
sine[3941] =70;
sine[3942] =70;
sine[3943] =70;
sine[3944] =70;
sine[3945] =69;
sine[3946] =69;
sine[3947] =69;
sine[3948] =69;
sine[3949] =68;
sine[3950] =68;
sine[3951] =68;
sine[3952] =68;
sine[3953] =67;
sine[3954] =67;
sine[3955] =67;
sine[3956] =66;
sine[3957] =66;
sine[3958] =66;
sine[3959] =66;
sine[3960] =65;
sine[3961] =65;
sine[3962] =65;
sine[3963] =65;
sine[3964] =64;
sine[3965] =64;
sine[3966] =64;
sine[3967] =64;
sine[3968] =63;
sine[3969] =63;
sine[3970] =63;
sine[3971] =63;
sine[3972] =62;
sine[3973] =62;
sine[3974] =62;
sine[3975] =62;
sine[3976] =61;
sine[3977] =61;
sine[3978] =61;
sine[3979] =61;
sine[3980] =60;
sine[3981] =60;
sine[3982] =60;
sine[3983] =59;
sine[3984] =59;
sine[3985] =59;
sine[3986] =59;
sine[3987] =58;
sine[3988] =58;
sine[3989] =58;
sine[3990] =58;
sine[3991] =57;
sine[3992] =57;
sine[3993] =57;
sine[3994] =57;
sine[3995] =57;
sine[3996] =56;
sine[3997] =56;
sine[3998] =56;
sine[3999] =56;
sine[4000] =55;
sine[4001] =55;
sine[4002] =55;
sine[4003] =55;
sine[4004] =54;
sine[4005] =54;
sine[4006] =54;
sine[4007] =54;
sine[4008] =53;
sine[4009] =53;
sine[4010] =53;
sine[4011] =53;
sine[4012] =52;
sine[4013] =52;
sine[4014] =52;
sine[4015] =52;
sine[4016] =51;
sine[4017] =51;
sine[4018] =51;
sine[4019] =51;
sine[4020] =51;
sine[4021] =50;
sine[4022] =50;
sine[4023] =50;
sine[4024] =50;
sine[4025] =49;
sine[4026] =49;
sine[4027] =49;
sine[4028] =49;
sine[4029] =48;
sine[4030] =48;
sine[4031] =48;
sine[4032] =48;
sine[4033] =48;
sine[4034] =47;
sine[4035] =47;
sine[4036] =47;
sine[4037] =47;
sine[4038] =46;
sine[4039] =46;
sine[4040] =46;
sine[4041] =46;
sine[4042] =45;
sine[4043] =45;
sine[4044] =45;
sine[4045] =45;
sine[4046] =45;
sine[4047] =44;
sine[4048] =44;
sine[4049] =44;
sine[4050] =44;
sine[4051] =43;
sine[4052] =43;
sine[4053] =43;
sine[4054] =43;
sine[4055] =43;
sine[4056] =42;
sine[4057] =42;
sine[4058] =42;
sine[4059] =42;
sine[4060] =42;
sine[4061] =41;
sine[4062] =41;
sine[4063] =41;
sine[4064] =41;
sine[4065] =40;
sine[4066] =40;
sine[4067] =40;
sine[4068] =40;
sine[4069] =40;
sine[4070] =39;
sine[4071] =39;
sine[4072] =39;
sine[4073] =39;
sine[4074] =39;
sine[4075] =38;
sine[4076] =38;
sine[4077] =38;
sine[4078] =38;
sine[4079] =38;
sine[4080] =37;
sine[4081] =37;
sine[4082] =37;
sine[4083] =37;
sine[4084] =37;
sine[4085] =36;
sine[4086] =36;
sine[4087] =36;
sine[4088] =36;
sine[4089] =36;
sine[4090] =35;
sine[4091] =35;
sine[4092] =35;
sine[4093] =35;
sine[4094] =35;
sine[4095] =34;
    end 
    
        always@ (posedge(Clk))
    begin
        data_out_3 = sine[k];
        k = k+ 1;
        if(k == 4095)
            k = 0;
    end
endmodule