module LUT_method_2(Clk,reset,data_out_2);
    input Clk,reset;
    output reg [11:0] data_out_2;
    reg [20:0] counter; 
    reg [11:0] sine [0:4095];
    integer j;  
    
    initial begin
        j = 0;
        sine[0] =477;
sine[1] =477;
sine[2] =476;
sine[3] =476;
sine[4] =476;
sine[5] =476;
sine[6] =476;
sine[7] =475;
sine[8] =475;
sine[9] =475;
sine[10] =475;
sine[11] =475;
sine[12] =474;
sine[13] =474;
sine[14] =474;
sine[15] =474;
sine[16] =474;
sine[17] =473;
sine[18] =473;
sine[19] =473;
sine[20] =473;
sine[21] =473;
sine[22] =472;
sine[23] =472;
sine[24] =472;
sine[25] =472;
sine[26] =472;
sine[27] =471;
sine[28] =471;
sine[29] =471;
sine[30] =471;
sine[31] =471;
sine[32] =470;
sine[33] =470;
sine[34] =470;
sine[35] =470;
sine[36] =469;
sine[37] =469;
sine[38] =469;
sine[39] =469;
sine[40] =469;
sine[41] =468;
sine[42] =468;
sine[43] =468;
sine[44] =468;
sine[45] =468;
sine[46] =467;
sine[47] =467;
sine[48] =467;
sine[49] =467;
sine[50] =466;
sine[51] =466;
sine[52] =466;
sine[53] =466;
sine[54] =466;
sine[55] =465;
sine[56] =465;
sine[57] =465;
sine[58] =465;
sine[59] =464;
sine[60] =464;
sine[61] =464;
sine[62] =464;
sine[63] =463;
sine[64] =463;
sine[65] =463;
sine[66] =463;
sine[67] =463;
sine[68] =462;
sine[69] =462;
sine[70] =462;
sine[71] =462;
sine[72] =461;
sine[73] =461;
sine[74] =461;
sine[75] =461;
sine[76] =460;
sine[77] =460;
sine[78] =460;
sine[79] =460;
sine[80] =460;
sine[81] =459;
sine[82] =459;
sine[83] =459;
sine[84] =459;
sine[85] =458;
sine[86] =458;
sine[87] =458;
sine[88] =458;
sine[89] =457;
sine[90] =457;
sine[91] =457;
sine[92] =457;
sine[93] =456;
sine[94] =456;
sine[95] =456;
sine[96] =456;
sine[97] =455;
sine[98] =455;
sine[99] =455;
sine[100] =455;
sine[101] =454;
sine[102] =454;
sine[103] =454;
sine[104] =454;
sine[105] =454;
sine[106] =453;
sine[107] =453;
sine[108] =453;
sine[109] =453;
sine[110] =452;
sine[111] =452;
sine[112] =452;
sine[113] =452;
sine[114] =451;
sine[115] =451;
sine[116] =451;
sine[117] =450;
sine[118] =450;
sine[119] =450;
sine[120] =450;
sine[121] =449;
sine[122] =449;
sine[123] =449;
sine[124] =449;
sine[125] =448;
sine[126] =448;
sine[127] =448;
sine[128] =448;
sine[129] =447;
sine[130] =447;
sine[131] =447;
sine[132] =447;
sine[133] =446;
sine[134] =446;
sine[135] =446;
sine[136] =446;
sine[137] =445;
sine[138] =445;
sine[139] =445;
sine[140] =445;
sine[141] =444;
sine[142] =444;
sine[143] =444;
sine[144] =443;
sine[145] =443;
sine[146] =443;
sine[147] =443;
sine[148] =442;
sine[149] =442;
sine[150] =442;
sine[151] =442;
sine[152] =441;
sine[153] =441;
sine[154] =441;
sine[155] =441;
sine[156] =440;
sine[157] =440;
sine[158] =440;
sine[159] =439;
sine[160] =439;
sine[161] =439;
sine[162] =439;
sine[163] =438;
sine[164] =438;
sine[165] =438;
sine[166] =438;
sine[167] =437;
sine[168] =437;
sine[169] =437;
sine[170] =436;
sine[171] =436;
sine[172] =436;
sine[173] =436;
sine[174] =435;
sine[175] =435;
sine[176] =435;
sine[177] =434;
sine[178] =434;
sine[179] =434;
sine[180] =434;
sine[181] =433;
sine[182] =433;
sine[183] =433;
sine[184] =433;
sine[185] =432;
sine[186] =432;
sine[187] =432;
sine[188] =431;
sine[189] =431;
sine[190] =431;
sine[191] =431;
sine[192] =430;
sine[193] =430;
sine[194] =430;
sine[195] =429;
sine[196] =429;
sine[197] =429;
sine[198] =429;
sine[199] =428;
sine[200] =428;
sine[201] =428;
sine[202] =427;
sine[203] =427;
sine[204] =427;
sine[205] =427;
sine[206] =426;
sine[207] =426;
sine[208] =426;
sine[209] =425;
sine[210] =425;
sine[211] =425;
sine[212] =424;
sine[213] =424;
sine[214] =424;
sine[215] =424;
sine[216] =423;
sine[217] =423;
sine[218] =423;
sine[219] =422;
sine[220] =422;
sine[221] =422;
sine[222] =421;
sine[223] =421;
sine[224] =421;
sine[225] =421;
sine[226] =420;
sine[227] =420;
sine[228] =420;
sine[229] =419;
sine[230] =419;
sine[231] =419;
sine[232] =418;
sine[233] =418;
sine[234] =418;
sine[235] =418;
sine[236] =417;
sine[237] =417;
sine[238] =417;
sine[239] =416;
sine[240] =416;
sine[241] =416;
sine[242] =415;
sine[243] =415;
sine[244] =415;
sine[245] =415;
sine[246] =414;
sine[247] =414;
sine[248] =414;
sine[249] =413;
sine[250] =413;
sine[251] =413;
sine[252] =412;
sine[253] =412;
sine[254] =412;
sine[255] =411;
sine[256] =411;
sine[257] =411;
sine[258] =411;
sine[259] =410;
sine[260] =410;
sine[261] =410;
sine[262] =409;
sine[263] =409;
sine[264] =409;
sine[265] =408;
sine[266] =408;
sine[267] =408;
sine[268] =407;
sine[269] =407;
sine[270] =407;
sine[271] =406;
sine[272] =406;
sine[273] =406;
sine[274] =405;
sine[275] =405;
sine[276] =405;
sine[277] =405;
sine[278] =404;
sine[279] =404;
sine[280] =404;
sine[281] =403;
sine[282] =403;
sine[283] =403;
sine[284] =402;
sine[285] =402;
sine[286] =402;
sine[287] =401;
sine[288] =401;
sine[289] =401;
sine[290] =400;
sine[291] =400;
sine[292] =400;
sine[293] =399;
sine[294] =399;
sine[295] =399;
sine[296] =398;
sine[297] =398;
sine[298] =398;
sine[299] =397;
sine[300] =397;
sine[301] =397;
sine[302] =396;
sine[303] =396;
sine[304] =396;
sine[305] =395;
sine[306] =395;
sine[307] =395;
sine[308] =395;
sine[309] =394;
sine[310] =394;
sine[311] =394;
sine[312] =393;
sine[313] =393;
sine[314] =393;
sine[315] =392;
sine[316] =392;
sine[317] =392;
sine[318] =391;
sine[319] =391;
sine[320] =391;
sine[321] =390;
sine[322] =390;
sine[323] =390;
sine[324] =389;
sine[325] =389;
sine[326] =389;
sine[327] =388;
sine[328] =388;
sine[329] =388;
sine[330] =387;
sine[331] =387;
sine[332] =387;
sine[333] =386;
sine[334] =386;
sine[335] =386;
sine[336] =385;
sine[337] =385;
sine[338] =384;
sine[339] =384;
sine[340] =384;
sine[341] =383;
sine[342] =383;
sine[343] =383;
sine[344] =382;
sine[345] =382;
sine[346] =382;
sine[347] =381;
sine[348] =381;
sine[349] =381;
sine[350] =380;
sine[351] =380;
sine[352] =380;
sine[353] =379;
sine[354] =379;
sine[355] =379;
sine[356] =378;
sine[357] =378;
sine[358] =378;
sine[359] =377;
sine[360] =377;
sine[361] =377;
sine[362] =376;
sine[363] =376;
sine[364] =376;
sine[365] =375;
sine[366] =375;
sine[367] =375;
sine[368] =374;
sine[369] =374;
sine[370] =374;
sine[371] =373;
sine[372] =373;
sine[373] =372;
sine[374] =372;
sine[375] =372;
sine[376] =371;
sine[377] =371;
sine[378] =371;
sine[379] =370;
sine[380] =370;
sine[381] =370;
sine[382] =369;
sine[383] =369;
sine[384] =369;
sine[385] =368;
sine[386] =368;
sine[387] =368;
sine[388] =367;
sine[389] =367;
sine[390] =367;
sine[391] =366;
sine[392] =366;
sine[393] =365;
sine[394] =365;
sine[395] =365;
sine[396] =364;
sine[397] =364;
sine[398] =364;
sine[399] =363;
sine[400] =363;
sine[401] =363;
sine[402] =362;
sine[403] =362;
sine[404] =362;
sine[405] =361;
sine[406] =361;
sine[407] =360;
sine[408] =360;
sine[409] =360;
sine[410] =359;
sine[411] =359;
sine[412] =359;
sine[413] =358;
sine[414] =358;
sine[415] =358;
sine[416] =357;
sine[417] =357;
sine[418] =357;
sine[419] =356;
sine[420] =356;
sine[421] =355;
sine[422] =355;
sine[423] =355;
sine[424] =354;
sine[425] =354;
sine[426] =354;
sine[427] =353;
sine[428] =353;
sine[429] =353;
sine[430] =352;
sine[431] =352;
sine[432] =351;
sine[433] =351;
sine[434] =351;
sine[435] =350;
sine[436] =350;
sine[437] =350;
sine[438] =349;
sine[439] =349;
sine[440] =349;
sine[441] =348;
sine[442] =348;
sine[443] =347;
sine[444] =347;
sine[445] =347;
sine[446] =346;
sine[447] =346;
sine[448] =346;
sine[449] =345;
sine[450] =345;
sine[451] =345;
sine[452] =344;
sine[453] =344;
sine[454] =343;
sine[455] =343;
sine[456] =343;
sine[457] =342;
sine[458] =342;
sine[459] =342;
sine[460] =341;
sine[461] =341;
sine[462] =340;
sine[463] =340;
sine[464] =340;
sine[465] =339;
sine[466] =339;
sine[467] =339;
sine[468] =338;
sine[469] =338;
sine[470] =338;
sine[471] =337;
sine[472] =337;
sine[473] =336;
sine[474] =336;
sine[475] =336;
sine[476] =335;
sine[477] =335;
sine[478] =335;
sine[479] =334;
sine[480] =334;
sine[481] =333;
sine[482] =333;
sine[483] =333;
sine[484] =332;
sine[485] =332;
sine[486] =332;
sine[487] =331;
sine[488] =331;
sine[489] =330;
sine[490] =330;
sine[491] =330;
sine[492] =329;
sine[493] =329;
sine[494] =329;
sine[495] =328;
sine[496] =328;
sine[497] =327;
sine[498] =327;
sine[499] =327;
sine[500] =326;
sine[501] =326;
sine[502] =326;
sine[503] =325;
sine[504] =325;
sine[505] =324;
sine[506] =324;
sine[507] =324;
sine[508] =323;
sine[509] =323;
sine[510] =323;
sine[511] =322;
sine[512] =322;
sine[513] =321;
sine[514] =321;
sine[515] =321;
sine[516] =320;
sine[517] =320;
sine[518] =319;
sine[519] =319;
sine[520] =319;
sine[521] =318;
sine[522] =318;
sine[523] =318;
sine[524] =317;
sine[525] =317;
sine[526] =316;
sine[527] =316;
sine[528] =316;
sine[529] =315;
sine[530] =315;
sine[531] =315;
sine[532] =314;
sine[533] =314;
sine[534] =313;
sine[535] =313;
sine[536] =313;
sine[537] =312;
sine[538] =312;
sine[539] =311;
sine[540] =311;
sine[541] =311;
sine[542] =310;
sine[543] =310;
sine[544] =310;
sine[545] =309;
sine[546] =309;
sine[547] =308;
sine[548] =308;
sine[549] =308;
sine[550] =307;
sine[551] =307;
sine[552] =306;
sine[553] =306;
sine[554] =306;
sine[555] =305;
sine[556] =305;
sine[557] =305;
sine[558] =304;
sine[559] =304;
sine[560] =303;
sine[561] =303;
sine[562] =303;
sine[563] =302;
sine[564] =302;
sine[565] =301;
sine[566] =301;
sine[567] =301;
sine[568] =300;
sine[569] =300;
sine[570] =300;
sine[571] =299;
sine[572] =299;
sine[573] =298;
sine[574] =298;
sine[575] =298;
sine[576] =297;
sine[577] =297;
sine[578] =296;
sine[579] =296;
sine[580] =296;
sine[581] =295;
sine[582] =295;
sine[583] =295;
sine[584] =294;
sine[585] =294;
sine[586] =293;
sine[587] =293;
sine[588] =293;
sine[589] =292;
sine[590] =292;
sine[591] =291;
sine[592] =291;
sine[593] =291;
sine[594] =290;
sine[595] =290;
sine[596] =289;
sine[597] =289;
sine[598] =289;
sine[599] =288;
sine[600] =288;
sine[601] =288;
sine[602] =287;
sine[603] =287;
sine[604] =286;
sine[605] =286;
sine[606] =286;
sine[607] =285;
sine[608] =285;
sine[609] =284;
sine[610] =284;
sine[611] =284;
sine[612] =283;
sine[613] =283;
sine[614] =282;
sine[615] =282;
sine[616] =282;
sine[617] =281;
sine[618] =281;
sine[619] =281;
sine[620] =280;
sine[621] =280;
sine[622] =279;
sine[623] =279;
sine[624] =279;
sine[625] =278;
sine[626] =278;
sine[627] =277;
sine[628] =277;
sine[629] =277;
sine[630] =276;
sine[631] =276;
sine[632] =275;
sine[633] =275;
sine[634] =275;
sine[635] =274;
sine[636] =274;
sine[637] =274;
sine[638] =273;
sine[639] =273;
sine[640] =272;
sine[641] =272;
sine[642] =272;
sine[643] =271;
sine[644] =271;
sine[645] =270;
sine[646] =270;
sine[647] =270;
sine[648] =269;
sine[649] =269;
sine[650] =268;
sine[651] =268;
sine[652] =268;
sine[653] =267;
sine[654] =267;
sine[655] =266;
sine[656] =266;
sine[657] =266;
sine[658] =265;
sine[659] =265;
sine[660] =265;
sine[661] =264;
sine[662] =264;
sine[663] =263;
sine[664] =263;
sine[665] =263;
sine[666] =262;
sine[667] =262;
sine[668] =261;
sine[669] =261;
sine[670] =261;
sine[671] =260;
sine[672] =260;
sine[673] =259;
sine[674] =259;
sine[675] =259;
sine[676] =258;
sine[677] =258;
sine[678] =257;
sine[679] =257;
sine[680] =257;
sine[681] =256;
sine[682] =256;
sine[683] =256;
sine[684] =255;
sine[685] =255;
sine[686] =254;
sine[687] =254;
sine[688] =254;
sine[689] =253;
sine[690] =253;
sine[691] =252;
sine[692] =252;
sine[693] =252;
sine[694] =251;
sine[695] =251;
sine[696] =250;
sine[697] =250;
sine[698] =250;
sine[699] =249;
sine[700] =249;
sine[701] =248;
sine[702] =248;
sine[703] =248;
sine[704] =247;
sine[705] =247;
sine[706] =246;
sine[707] =246;
sine[708] =246;
sine[709] =245;
sine[710] =245;
sine[711] =245;
sine[712] =244;
sine[713] =244;
sine[714] =243;
sine[715] =243;
sine[716] =243;
sine[717] =242;
sine[718] =242;
sine[719] =241;
sine[720] =241;
sine[721] =241;
sine[722] =240;
sine[723] =240;
sine[724] =239;
sine[725] =239;
sine[726] =239;
sine[727] =238;
sine[728] =238;
sine[729] =237;
sine[730] =237;
sine[731] =237;
sine[732] =236;
sine[733] =236;
sine[734] =236;
sine[735] =235;
sine[736] =235;
sine[737] =234;
sine[738] =234;
sine[739] =234;
sine[740] =233;
sine[741] =233;
sine[742] =232;
sine[743] =232;
sine[744] =232;
sine[745] =231;
sine[746] =231;
sine[747] =230;
sine[748] =230;
sine[749] =230;
sine[750] =229;
sine[751] =229;
sine[752] =229;
sine[753] =228;
sine[754] =228;
sine[755] =227;
sine[756] =227;
sine[757] =227;
sine[758] =226;
sine[759] =226;
sine[760] =225;
sine[761] =225;
sine[762] =225;
sine[763] =224;
sine[764] =224;
sine[765] =223;
sine[766] =223;
sine[767] =223;
sine[768] =222;
sine[769] =222;
sine[770] =222;
sine[771] =221;
sine[772] =221;
sine[773] =220;
sine[774] =220;
sine[775] =220;
sine[776] =219;
sine[777] =219;
sine[778] =218;
sine[779] =218;
sine[780] =218;
sine[781] =217;
sine[782] =217;
sine[783] =216;
sine[784] =216;
sine[785] =216;
sine[786] =215;
sine[787] =215;
sine[788] =215;
sine[789] =214;
sine[790] =214;
sine[791] =213;
sine[792] =213;
sine[793] =213;
sine[794] =212;
sine[795] =212;
sine[796] =211;
sine[797] =211;
sine[798] =211;
sine[799] =210;
sine[800] =210;
sine[801] =210;
sine[802] =209;
sine[803] =209;
sine[804] =208;
sine[805] =208;
sine[806] =208;
sine[807] =207;
sine[808] =207;
sine[809] =206;
sine[810] =206;
sine[811] =206;
sine[812] =205;
sine[813] =205;
sine[814] =205;
sine[815] =204;
sine[816] =204;
sine[817] =203;
sine[818] =203;
sine[819] =203;
sine[820] =202;
sine[821] =202;
sine[822] =201;
sine[823] =201;
sine[824] =201;
sine[825] =200;
sine[826] =200;
sine[827] =200;
sine[828] =199;
sine[829] =199;
sine[830] =198;
sine[831] =198;
sine[832] =198;
sine[833] =197;
sine[834] =197;
sine[835] =196;
sine[836] =196;
sine[837] =196;
sine[838] =195;
sine[839] =195;
sine[840] =195;
sine[841] =194;
sine[842] =194;
sine[843] =193;
sine[844] =193;
sine[845] =193;
sine[846] =192;
sine[847] =192;
sine[848] =192;
sine[849] =191;
sine[850] =191;
sine[851] =190;
sine[852] =190;
sine[853] =190;
sine[854] =189;
sine[855] =189;
sine[856] =188;
sine[857] =188;
sine[858] =188;
sine[859] =187;
sine[860] =187;
sine[861] =187;
sine[862] =186;
sine[863] =186;
sine[864] =185;
sine[865] =185;
sine[866] =185;
sine[867] =184;
sine[868] =184;
sine[869] =184;
sine[870] =183;
sine[871] =183;
sine[872] =182;
sine[873] =182;
sine[874] =182;
sine[875] =181;
sine[876] =181;
sine[877] =181;
sine[878] =180;
sine[879] =180;
sine[880] =179;
sine[881] =179;
sine[882] =179;
sine[883] =178;
sine[884] =178;
sine[885] =178;
sine[886] =177;
sine[887] =177;
sine[888] =176;
sine[889] =176;
sine[890] =176;
sine[891] =175;
sine[892] =175;
sine[893] =175;
sine[894] =174;
sine[895] =174;
sine[896] =173;
sine[897] =173;
sine[898] =173;
sine[899] =172;
sine[900] =172;
sine[901] =172;
sine[902] =171;
sine[903] =171;
sine[904] =171;
sine[905] =170;
sine[906] =170;
sine[907] =169;
sine[908] =169;
sine[909] =169;
sine[910] =168;
sine[911] =168;
sine[912] =168;
sine[913] =167;
sine[914] =167;
sine[915] =166;
sine[916] =166;
sine[917] =166;
sine[918] =165;
sine[919] =165;
sine[920] =165;
sine[921] =164;
sine[922] =164;
sine[923] =164;
sine[924] =163;
sine[925] =163;
sine[926] =162;
sine[927] =162;
sine[928] =162;
sine[929] =161;
sine[930] =161;
sine[931] =161;
sine[932] =160;
sine[933] =160;
sine[934] =160;
sine[935] =159;
sine[936] =159;
sine[937] =158;
sine[938] =158;
sine[939] =158;
sine[940] =157;
sine[941] =157;
sine[942] =157;
sine[943] =156;
sine[944] =156;
sine[945] =156;
sine[946] =155;
sine[947] =155;
sine[948] =154;
sine[949] =154;
sine[950] =154;
sine[951] =153;
sine[952] =153;
sine[953] =153;
sine[954] =152;
sine[955] =152;
sine[956] =152;
sine[957] =151;
sine[958] =151;
sine[959] =151;
sine[960] =150;
sine[961] =150;
sine[962] =149;
sine[963] =149;
sine[964] =149;
sine[965] =148;
sine[966] =148;
sine[967] =148;
sine[968] =147;
sine[969] =147;
sine[970] =147;
sine[971] =146;
sine[972] =146;
sine[973] =146;
sine[974] =145;
sine[975] =145;
sine[976] =144;
sine[977] =144;
sine[978] =144;
sine[979] =143;
sine[980] =143;
sine[981] =143;
sine[982] =142;
sine[983] =142;
sine[984] =142;
sine[985] =141;
sine[986] =141;
sine[987] =141;
sine[988] =140;
sine[989] =140;
sine[990] =140;
sine[991] =139;
sine[992] =139;
sine[993] =139;
sine[994] =138;
sine[995] =138;
sine[996] =137;
sine[997] =137;
sine[998] =137;
sine[999] =136;
sine[1000] =136;
sine[1001] =136;
sine[1002] =135;
sine[1003] =135;
sine[1004] =135;
sine[1005] =134;
sine[1006] =134;
sine[1007] =134;
sine[1008] =133;
sine[1009] =133;
sine[1010] =133;
sine[1011] =132;
sine[1012] =132;
sine[1013] =132;
sine[1014] =131;
sine[1015] =131;
sine[1016] =131;
sine[1017] =130;
sine[1018] =130;
sine[1019] =130;
sine[1020] =129;
sine[1021] =129;
sine[1022] =129;
sine[1023] =128;
sine[1024] =128;
sine[1025] =128;
sine[1026] =127;
sine[1027] =127;
sine[1028] =127;
sine[1029] =126;
sine[1030] =126;
sine[1031] =125;
sine[1032] =125;
sine[1033] =125;
sine[1034] =124;
sine[1035] =124;
sine[1036] =124;
sine[1037] =123;
sine[1038] =123;
sine[1039] =123;
sine[1040] =122;
sine[1041] =122;
sine[1042] =122;
sine[1043] =121;
sine[1044] =121;
sine[1045] =121;
sine[1046] =120;
sine[1047] =120;
sine[1048] =120;
sine[1049] =119;
sine[1050] =119;
sine[1051] =119;
sine[1052] =118;
sine[1053] =118;
sine[1054] =118;
sine[1055] =117;
sine[1056] =117;
sine[1057] =117;
sine[1058] =116;
sine[1059] =116;
sine[1060] =116;
sine[1061] =116;
sine[1062] =115;
sine[1063] =115;
sine[1064] =115;
sine[1065] =114;
sine[1066] =114;
sine[1067] =114;
sine[1068] =113;
sine[1069] =113;
sine[1070] =113;
sine[1071] =112;
sine[1072] =112;
sine[1073] =112;
sine[1074] =111;
sine[1075] =111;
sine[1076] =111;
sine[1077] =110;
sine[1078] =110;
sine[1079] =110;
sine[1080] =109;
sine[1081] =109;
sine[1082] =109;
sine[1083] =108;
sine[1084] =108;
sine[1085] =108;
sine[1086] =107;
sine[1087] =107;
sine[1088] =107;
sine[1089] =106;
sine[1090] =106;
sine[1091] =106;
sine[1092] =106;
sine[1093] =105;
sine[1094] =105;
sine[1095] =105;
sine[1096] =104;
sine[1097] =104;
sine[1098] =104;
sine[1099] =103;
sine[1100] =103;
sine[1101] =103;
sine[1102] =102;
sine[1103] =102;
sine[1104] =102;
sine[1105] =101;
sine[1106] =101;
sine[1107] =101;
sine[1108] =100;
sine[1109] =100;
sine[1110] =100;
sine[1111] =100;
sine[1112] =99;
sine[1113] =99;
sine[1114] =99;
sine[1115] =98;
sine[1116] =98;
sine[1117] =98;
sine[1118] =97;
sine[1119] =97;
sine[1120] =97;
sine[1121] =96;
sine[1122] =96;
sine[1123] =96;
sine[1124] =96;
sine[1125] =95;
sine[1126] =95;
sine[1127] =95;
sine[1128] =94;
sine[1129] =94;
sine[1130] =94;
sine[1131] =93;
sine[1132] =93;
sine[1133] =93;
sine[1134] =93;
sine[1135] =92;
sine[1136] =92;
sine[1137] =92;
sine[1138] =91;
sine[1139] =91;
sine[1140] =91;
sine[1141] =90;
sine[1142] =90;
sine[1143] =90;
sine[1144] =90;
sine[1145] =89;
sine[1146] =89;
sine[1147] =89;
sine[1148] =88;
sine[1149] =88;
sine[1150] =88;
sine[1151] =87;
sine[1152] =87;
sine[1153] =87;
sine[1154] =87;
sine[1155] =86;
sine[1156] =86;
sine[1157] =86;
sine[1158] =85;
sine[1159] =85;
sine[1160] =85;
sine[1161] =84;
sine[1162] =84;
sine[1163] =84;
sine[1164] =84;
sine[1165] =83;
sine[1166] =83;
sine[1167] =83;
sine[1168] =82;
sine[1169] =82;
sine[1170] =82;
sine[1171] =82;
sine[1172] =81;
sine[1173] =81;
sine[1174] =81;
sine[1175] =80;
sine[1176] =80;
sine[1177] =80;
sine[1178] =80;
sine[1179] =79;
sine[1180] =79;
sine[1181] =79;
sine[1182] =78;
sine[1183] =78;
sine[1184] =78;
sine[1185] =78;
sine[1186] =77;
sine[1187] =77;
sine[1188] =77;
sine[1189] =77;
sine[1190] =76;
sine[1191] =76;
sine[1192] =76;
sine[1193] =75;
sine[1194] =75;
sine[1195] =75;
sine[1196] =75;
sine[1197] =74;
sine[1198] =74;
sine[1199] =74;
sine[1200] =73;
sine[1201] =73;
sine[1202] =73;
sine[1203] =73;
sine[1204] =72;
sine[1205] =72;
sine[1206] =72;
sine[1207] =72;
sine[1208] =71;
sine[1209] =71;
sine[1210] =71;
sine[1211] =70;
sine[1212] =70;
sine[1213] =70;
sine[1214] =70;
sine[1215] =69;
sine[1216] =69;
sine[1217] =69;
sine[1218] =69;
sine[1219] =68;
sine[1220] =68;
sine[1221] =68;
sine[1222] =68;
sine[1223] =67;
sine[1224] =67;
sine[1225] =67;
sine[1226] =66;
sine[1227] =66;
sine[1228] =66;
sine[1229] =66;
sine[1230] =65;
sine[1231] =65;
sine[1232] =65;
sine[1233] =65;
sine[1234] =64;
sine[1235] =64;
sine[1236] =64;
sine[1237] =64;
sine[1238] =63;
sine[1239] =63;
sine[1240] =63;
sine[1241] =63;
sine[1242] =62;
sine[1243] =62;
sine[1244] =62;
sine[1245] =62;
sine[1246] =61;
sine[1247] =61;
sine[1248] =61;
sine[1249] =61;
sine[1250] =60;
sine[1251] =60;
sine[1252] =60;
sine[1253] =59;
sine[1254] =59;
sine[1255] =59;
sine[1256] =59;
sine[1257] =58;
sine[1258] =58;
sine[1259] =58;
sine[1260] =58;
sine[1261] =57;
sine[1262] =57;
sine[1263] =57;
sine[1264] =57;
sine[1265] =57;
sine[1266] =56;
sine[1267] =56;
sine[1268] =56;
sine[1269] =56;
sine[1270] =55;
sine[1271] =55;
sine[1272] =55;
sine[1273] =55;
sine[1274] =54;
sine[1275] =54;
sine[1276] =54;
sine[1277] =54;
sine[1278] =53;
sine[1279] =53;
sine[1280] =53;
sine[1281] =53;
sine[1282] =52;
sine[1283] =52;
sine[1284] =52;
sine[1285] =52;
sine[1286] =51;
sine[1287] =51;
sine[1288] =51;
sine[1289] =51;
sine[1290] =51;
sine[1291] =50;
sine[1292] =50;
sine[1293] =50;
sine[1294] =50;
sine[1295] =49;
sine[1296] =49;
sine[1297] =49;
sine[1298] =49;
sine[1299] =48;
sine[1300] =48;
sine[1301] =48;
sine[1302] =48;
sine[1303] =48;
sine[1304] =47;
sine[1305] =47;
sine[1306] =47;
sine[1307] =47;
sine[1308] =46;
sine[1309] =46;
sine[1310] =46;
sine[1311] =46;
sine[1312] =45;
sine[1313] =45;
sine[1314] =45;
sine[1315] =45;
sine[1316] =45;
sine[1317] =44;
sine[1318] =44;
sine[1319] =44;
sine[1320] =44;
sine[1321] =43;
sine[1322] =43;
sine[1323] =43;
sine[1324] =43;
sine[1325] =43;
sine[1326] =42;
sine[1327] =42;
sine[1328] =42;
sine[1329] =42;
sine[1330] =42;
sine[1331] =41;
sine[1332] =41;
sine[1333] =41;
sine[1334] =41;
sine[1335] =40;
sine[1336] =40;
sine[1337] =40;
sine[1338] =40;
sine[1339] =40;
sine[1340] =39;
sine[1341] =39;
sine[1342] =39;
sine[1343] =39;
sine[1344] =39;
sine[1345] =38;
sine[1346] =38;
sine[1347] =38;
sine[1348] =38;
sine[1349] =38;
sine[1350] =37;
sine[1351] =37;
sine[1352] =37;
sine[1353] =37;
sine[1354] =37;
sine[1355] =36;
sine[1356] =36;
sine[1357] =36;
sine[1358] =36;
sine[1359] =36;
sine[1360] =35;
sine[1361] =35;
sine[1362] =35;
sine[1363] =35;
sine[1364] =35;
sine[1365] =34;
sine[1366] =34;
sine[1367] =34;
sine[1368] =34;
sine[1369] =34;
sine[1370] =33;
sine[1371] =33;
sine[1372] =33;
sine[1373] =33;
sine[1374] =33;
sine[1375] =32;
sine[1376] =32;
sine[1377] =32;
sine[1378] =32;
sine[1379] =32;
sine[1380] =31;
sine[1381] =31;
sine[1382] =31;
sine[1383] =31;
sine[1384] =31;
sine[1385] =31;
sine[1386] =30;
sine[1387] =30;
sine[1388] =30;
sine[1389] =30;
sine[1390] =30;
sine[1391] =29;
sine[1392] =29;
sine[1393] =29;
sine[1394] =29;
sine[1395] =29;
sine[1396] =29;
sine[1397] =28;
sine[1398] =28;
sine[1399] =28;
sine[1400] =28;
sine[1401] =28;
sine[1402] =27;
sine[1403] =27;
sine[1404] =27;
sine[1405] =27;
sine[1406] =27;
sine[1407] =27;
sine[1408] =26;
sine[1409] =26;
sine[1410] =26;
sine[1411] =26;
sine[1412] =26;
sine[1413] =26;
sine[1414] =25;
sine[1415] =25;
sine[1416] =25;
sine[1417] =25;
sine[1418] =25;
sine[1419] =25;
sine[1420] =24;
sine[1421] =24;
sine[1422] =24;
sine[1423] =24;
sine[1424] =24;
sine[1425] =24;
sine[1426] =23;
sine[1427] =23;
sine[1428] =23;
sine[1429] =23;
sine[1430] =23;
sine[1431] =23;
sine[1432] =22;
sine[1433] =22;
sine[1434] =22;
sine[1435] =22;
sine[1436] =22;
sine[1437] =22;
sine[1438] =21;
sine[1439] =21;
sine[1440] =21;
sine[1441] =21;
sine[1442] =21;
sine[1443] =21;
sine[1444] =21;
sine[1445] =20;
sine[1446] =20;
sine[1447] =20;
sine[1448] =20;
sine[1449] =20;
sine[1450] =20;
sine[1451] =19;
sine[1452] =19;
sine[1453] =19;
sine[1454] =19;
sine[1455] =19;
sine[1456] =19;
sine[1457] =19;
sine[1458] =18;
sine[1459] =18;
sine[1460] =18;
sine[1461] =18;
sine[1462] =18;
sine[1463] =18;
sine[1464] =18;
sine[1465] =17;
sine[1466] =17;
sine[1467] =17;
sine[1468] =17;
sine[1469] =17;
sine[1470] =17;
sine[1471] =17;
sine[1472] =16;
sine[1473] =16;
sine[1474] =16;
sine[1475] =16;
sine[1476] =16;
sine[1477] =16;
sine[1478] =16;
sine[1479] =15;
sine[1480] =15;
sine[1481] =15;
sine[1482] =15;
sine[1483] =15;
sine[1484] =15;
sine[1485] =15;
sine[1486] =15;
sine[1487] =14;
sine[1488] =14;
sine[1489] =14;
sine[1490] =14;
sine[1491] =14;
sine[1492] =14;
sine[1493] =14;
sine[1494] =14;
sine[1495] =13;
sine[1496] =13;
sine[1497] =13;
sine[1498] =13;
sine[1499] =13;
sine[1500] =13;
sine[1501] =13;
sine[1502] =13;
sine[1503] =12;
sine[1504] =12;
sine[1505] =12;
sine[1506] =12;
sine[1507] =12;
sine[1508] =12;
sine[1509] =12;
sine[1510] =12;
sine[1511] =11;
sine[1512] =11;
sine[1513] =11;
sine[1514] =11;
sine[1515] =11;
sine[1516] =11;
sine[1517] =11;
sine[1518] =11;
sine[1519] =11;
sine[1520] =10;
sine[1521] =10;
sine[1522] =10;
sine[1523] =10;
sine[1524] =10;
sine[1525] =10;
sine[1526] =10;
sine[1527] =10;
sine[1528] =10;
sine[1529] =9;
sine[1530] =9;
sine[1531] =9;
sine[1532] =9;
sine[1533] =9;
sine[1534] =9;
sine[1535] =9;
sine[1536] =9;
sine[1537] =9;
sine[1538] =9;
sine[1539] =8;
sine[1540] =8;
sine[1541] =8;
sine[1542] =8;
sine[1543] =8;
sine[1544] =8;
sine[1545] =8;
sine[1546] =8;
sine[1547] =8;
sine[1548] =8;
sine[1549] =7;
sine[1550] =7;
sine[1551] =7;
sine[1552] =7;
sine[1553] =7;
sine[1554] =7;
sine[1555] =7;
sine[1556] =7;
sine[1557] =7;
sine[1558] =7;
sine[1559] =7;
sine[1560] =6;
sine[1561] =6;
sine[1562] =6;
sine[1563] =6;
sine[1564] =6;
sine[1565] =6;
sine[1566] =6;
sine[1567] =6;
sine[1568] =6;
sine[1569] =6;
sine[1570] =6;
sine[1571] =6;
sine[1572] =5;
sine[1573] =5;
sine[1574] =5;
sine[1575] =5;
sine[1576] =5;
sine[1577] =5;
sine[1578] =5;
sine[1579] =5;
sine[1580] =5;
sine[1581] =5;
sine[1582] =5;
sine[1583] =5;
sine[1584] =5;
sine[1585] =4;
sine[1586] =4;
sine[1587] =4;
sine[1588] =4;
sine[1589] =4;
sine[1590] =4;
sine[1591] =4;
sine[1592] =4;
sine[1593] =4;
sine[1594] =4;
sine[1595] =4;
sine[1596] =4;
sine[1597] =4;
sine[1598] =4;
sine[1599] =3;
sine[1600] =3;
sine[1601] =3;
sine[1602] =3;
sine[1603] =3;
sine[1604] =3;
sine[1605] =3;
sine[1606] =3;
sine[1607] =3;
sine[1608] =3;
sine[1609] =3;
sine[1610] =3;
sine[1611] =3;
sine[1612] =3;
sine[1613] =3;
sine[1614] =3;
sine[1615] =3;
sine[1616] =2;
sine[1617] =2;
sine[1618] =2;
sine[1619] =2;
sine[1620] =2;
sine[1621] =2;
sine[1622] =2;
sine[1623] =2;
sine[1624] =2;
sine[1625] =2;
sine[1626] =2;
sine[1627] =2;
sine[1628] =2;
sine[1629] =2;
sine[1630] =2;
sine[1631] =2;
sine[1632] =2;
sine[1633] =2;
sine[1634] =2;
sine[1635] =2;
sine[1636] =2;
sine[1637] =1;
sine[1638] =1;
sine[1639] =1;
sine[1640] =1;
sine[1641] =1;
sine[1642] =1;
sine[1643] =1;
sine[1644] =1;
sine[1645] =1;
sine[1646] =1;
sine[1647] =1;
sine[1648] =1;
sine[1649] =1;
sine[1650] =1;
sine[1651] =1;
sine[1652] =1;
sine[1653] =1;
sine[1654] =1;
sine[1655] =1;
sine[1656] =1;
sine[1657] =1;
sine[1658] =1;
sine[1659] =1;
sine[1660] =1;
sine[1661] =1;
sine[1662] =1;
sine[1663] =1;
sine[1664] =1;
sine[1665] =1;
sine[1666] =1;
sine[1667] =0;
sine[1668] =0;
sine[1669] =0;
sine[1670] =0;
sine[1671] =0;
sine[1672] =0;
sine[1673] =0;
sine[1674] =0;
sine[1675] =0;
sine[1676] =0;
sine[1677] =0;
sine[1678] =0;
sine[1679] =0;
sine[1680] =0;
sine[1681] =0;
sine[1682] =0;
sine[1683] =0;
sine[1684] =0;
sine[1685] =0;
sine[1686] =0;
sine[1687] =0;
sine[1688] =0;
sine[1689] =0;
sine[1690] =0;
sine[1691] =0;
sine[1692] =0;
sine[1693] =0;
sine[1694] =0;
sine[1695] =0;
sine[1696] =0;
sine[1697] =0;
sine[1698] =0;
sine[1699] =0;
sine[1700] =0;
sine[1701] =0;
sine[1702] =0;
sine[1703] =0;
sine[1704] =0;
sine[1705] =0;
sine[1706] =0;
sine[1707] =0;
sine[1708] =0;
sine[1709] =0;
sine[1710] =0;
sine[1711] =0;
sine[1712] =0;
sine[1713] =0;
sine[1714] =0;
sine[1715] =0;
sine[1716] =0;
sine[1717] =0;
sine[1718] =0;
sine[1719] =0;
sine[1720] =0;
sine[1721] =0;
sine[1722] =0;
sine[1723] =0;
sine[1724] =0;
sine[1725] =0;
sine[1726] =0;
sine[1727] =0;
sine[1728] =0;
sine[1729] =0;
sine[1730] =0;
sine[1731] =0;
sine[1732] =0;
sine[1733] =0;
sine[1734] =0;
sine[1735] =0;
sine[1736] =0;
sine[1737] =0;
sine[1738] =0;
sine[1739] =0;
sine[1740] =0;
sine[1741] =0;
sine[1742] =0;
sine[1743] =0;
sine[1744] =0;
sine[1745] =0;
sine[1746] =0;
sine[1747] =0;
sine[1748] =1;
sine[1749] =1;
sine[1750] =1;
sine[1751] =1;
sine[1752] =1;
sine[1753] =1;
sine[1754] =1;
sine[1755] =1;
sine[1756] =1;
sine[1757] =1;
sine[1758] =1;
sine[1759] =1;
sine[1760] =1;
sine[1761] =1;
sine[1762] =1;
sine[1763] =1;
sine[1764] =1;
sine[1765] =1;
sine[1766] =1;
sine[1767] =1;
sine[1768] =1;
sine[1769] =1;
sine[1770] =1;
sine[1771] =1;
sine[1772] =1;
sine[1773] =1;
sine[1774] =1;
sine[1775] =1;
sine[1776] =1;
sine[1777] =1;
sine[1778] =2;
sine[1779] =2;
sine[1780] =2;
sine[1781] =2;
sine[1782] =2;
sine[1783] =2;
sine[1784] =2;
sine[1785] =2;
sine[1786] =2;
sine[1787] =2;
sine[1788] =2;
sine[1789] =2;
sine[1790] =2;
sine[1791] =2;
sine[1792] =2;
sine[1793] =2;
sine[1794] =2;
sine[1795] =2;
sine[1796] =2;
sine[1797] =2;
sine[1798] =2;
sine[1799] =3;
sine[1800] =3;
sine[1801] =3;
sine[1802] =3;
sine[1803] =3;
sine[1804] =3;
sine[1805] =3;
sine[1806] =3;
sine[1807] =3;
sine[1808] =3;
sine[1809] =3;
sine[1810] =3;
sine[1811] =3;
sine[1812] =3;
sine[1813] =3;
sine[1814] =3;
sine[1815] =3;
sine[1816] =4;
sine[1817] =4;
sine[1818] =4;
sine[1819] =4;
sine[1820] =4;
sine[1821] =4;
sine[1822] =4;
sine[1823] =4;
sine[1824] =4;
sine[1825] =4;
sine[1826] =4;
sine[1827] =4;
sine[1828] =4;
sine[1829] =4;
sine[1830] =5;
sine[1831] =5;
sine[1832] =5;
sine[1833] =5;
sine[1834] =5;
sine[1835] =5;
sine[1836] =5;
sine[1837] =5;
sine[1838] =5;
sine[1839] =5;
sine[1840] =5;
sine[1841] =5;
sine[1842] =5;
sine[1843] =6;
sine[1844] =6;
sine[1845] =6;
sine[1846] =6;
sine[1847] =6;
sine[1848] =6;
sine[1849] =6;
sine[1850] =6;
sine[1851] =6;
sine[1852] =6;
sine[1853] =6;
sine[1854] =6;
sine[1855] =7;
sine[1856] =7;
sine[1857] =7;
sine[1858] =7;
sine[1859] =7;
sine[1860] =7;
sine[1861] =7;
sine[1862] =7;
sine[1863] =7;
sine[1864] =7;
sine[1865] =7;
sine[1866] =8;
sine[1867] =8;
sine[1868] =8;
sine[1869] =8;
sine[1870] =8;
sine[1871] =8;
sine[1872] =8;
sine[1873] =8;
sine[1874] =8;
sine[1875] =8;
sine[1876] =9;
sine[1877] =9;
sine[1878] =9;
sine[1879] =9;
sine[1880] =9;
sine[1881] =9;
sine[1882] =9;
sine[1883] =9;
sine[1884] =9;
sine[1885] =9;
sine[1886] =10;
sine[1887] =10;
sine[1888] =10;
sine[1889] =10;
sine[1890] =10;
sine[1891] =10;
sine[1892] =10;
sine[1893] =10;
sine[1894] =10;
sine[1895] =11;
sine[1896] =11;
sine[1897] =11;
sine[1898] =11;
sine[1899] =11;
sine[1900] =11;
sine[1901] =11;
sine[1902] =11;
sine[1903] =11;
sine[1904] =12;
sine[1905] =12;
sine[1906] =12;
sine[1907] =12;
sine[1908] =12;
sine[1909] =12;
sine[1910] =12;
sine[1911] =12;
sine[1912] =13;
sine[1913] =13;
sine[1914] =13;
sine[1915] =13;
sine[1916] =13;
sine[1917] =13;
sine[1918] =13;
sine[1919] =13;
sine[1920] =14;
sine[1921] =14;
sine[1922] =14;
sine[1923] =14;
sine[1924] =14;
sine[1925] =14;
sine[1926] =14;
sine[1927] =14;
sine[1928] =15;
sine[1929] =15;
sine[1930] =15;
sine[1931] =15;
sine[1932] =15;
sine[1933] =15;
sine[1934] =15;
sine[1935] =15;
sine[1936] =16;
sine[1937] =16;
sine[1938] =16;
sine[1939] =16;
sine[1940] =16;
sine[1941] =16;
sine[1942] =16;
sine[1943] =17;
sine[1944] =17;
sine[1945] =17;
sine[1946] =17;
sine[1947] =17;
sine[1948] =17;
sine[1949] =17;
sine[1950] =18;
sine[1951] =18;
sine[1952] =18;
sine[1953] =18;
sine[1954] =18;
sine[1955] =18;
sine[1956] =18;
sine[1957] =19;
sine[1958] =19;
sine[1959] =19;
sine[1960] =19;
sine[1961] =19;
sine[1962] =19;
sine[1963] =19;
sine[1964] =20;
sine[1965] =20;
sine[1966] =20;
sine[1967] =20;
sine[1968] =20;
sine[1969] =20;
sine[1970] =21;
sine[1971] =21;
sine[1972] =21;
sine[1973] =21;
sine[1974] =21;
sine[1975] =21;
sine[1976] =21;
sine[1977] =22;
sine[1978] =22;
sine[1979] =22;
sine[1980] =22;
sine[1981] =22;
sine[1982] =22;
sine[1983] =23;
sine[1984] =23;
sine[1985] =23;
sine[1986] =23;
sine[1987] =23;
sine[1988] =23;
sine[1989] =24;
sine[1990] =24;
sine[1991] =24;
sine[1992] =24;
sine[1993] =24;
sine[1994] =24;
sine[1995] =25;
sine[1996] =25;
sine[1997] =25;
sine[1998] =25;
sine[1999] =25;
sine[2000] =25;
sine[2001] =26;
sine[2002] =26;
sine[2003] =26;
sine[2004] =26;
sine[2005] =26;
sine[2006] =26;
sine[2007] =27;
sine[2008] =27;
sine[2009] =27;
sine[2010] =27;
sine[2011] =27;
sine[2012] =27;
sine[2013] =28;
sine[2014] =28;
sine[2015] =28;
sine[2016] =28;
sine[2017] =28;
sine[2018] =29;
sine[2019] =29;
sine[2020] =29;
sine[2021] =29;
sine[2022] =29;
sine[2023] =29;
sine[2024] =30;
sine[2025] =30;
sine[2026] =30;
sine[2027] =30;
sine[2028] =30;
sine[2029] =31;
sine[2030] =31;
sine[2031] =31;
sine[2032] =31;
sine[2033] =31;
sine[2034] =31;
sine[2035] =32;
sine[2036] =32;
sine[2037] =32;
sine[2038] =32;
sine[2039] =32;
sine[2040] =33;
sine[2041] =33;
sine[2042] =33;
sine[2043] =33;
sine[2044] =33;
sine[2045] =34;
sine[2046] =34;
sine[2047] =34;
sine[2048] =34;
sine[2049] =34;
sine[2050] =35;
sine[2051] =35;
sine[2052] =35;
sine[2053] =35;
sine[2054] =35;
sine[2055] =36;
sine[2056] =36;
sine[2057] =36;
sine[2058] =36;
sine[2059] =36;
sine[2060] =37;
sine[2061] =37;
sine[2062] =37;
sine[2063] =37;
sine[2064] =37;
sine[2065] =38;
sine[2066] =38;
sine[2067] =38;
sine[2068] =38;
sine[2069] =38;
sine[2070] =39;
sine[2071] =39;
sine[2072] =39;
sine[2073] =39;
sine[2074] =39;
sine[2075] =40;
sine[2076] =40;
sine[2077] =40;
sine[2078] =40;
sine[2079] =40;
sine[2080] =41;
sine[2081] =41;
sine[2082] =41;
sine[2083] =41;
sine[2084] =42;
sine[2085] =42;
sine[2086] =42;
sine[2087] =42;
sine[2088] =42;
sine[2089] =43;
sine[2090] =43;
sine[2091] =43;
sine[2092] =43;
sine[2093] =43;
sine[2094] =44;
sine[2095] =44;
sine[2096] =44;
sine[2097] =44;
sine[2098] =45;
sine[2099] =45;
sine[2100] =45;
sine[2101] =45;
sine[2102] =45;
sine[2103] =46;
sine[2104] =46;
sine[2105] =46;
sine[2106] =46;
sine[2107] =47;
sine[2108] =47;
sine[2109] =47;
sine[2110] =47;
sine[2111] =48;
sine[2112] =48;
sine[2113] =48;
sine[2114] =48;
sine[2115] =48;
sine[2116] =49;
sine[2117] =49;
sine[2118] =49;
sine[2119] =49;
sine[2120] =50;
sine[2121] =50;
sine[2122] =50;
sine[2123] =50;
sine[2124] =51;
sine[2125] =51;
sine[2126] =51;
sine[2127] =51;
sine[2128] =51;
sine[2129] =52;
sine[2130] =52;
sine[2131] =52;
sine[2132] =52;
sine[2133] =53;
sine[2134] =53;
sine[2135] =53;
sine[2136] =53;
sine[2137] =54;
sine[2138] =54;
sine[2139] =54;
sine[2140] =54;
sine[2141] =55;
sine[2142] =55;
sine[2143] =55;
sine[2144] =55;
sine[2145] =56;
sine[2146] =56;
sine[2147] =56;
sine[2148] =56;
sine[2149] =57;
sine[2150] =57;
sine[2151] =57;
sine[2152] =57;
sine[2153] =57;
sine[2154] =58;
sine[2155] =58;
sine[2156] =58;
sine[2157] =58;
sine[2158] =59;
sine[2159] =59;
sine[2160] =59;
sine[2161] =59;
sine[2162] =60;
sine[2163] =60;
sine[2164] =60;
sine[2165] =61;
sine[2166] =61;
sine[2167] =61;
sine[2168] =61;
sine[2169] =62;
sine[2170] =62;
sine[2171] =62;
sine[2172] =62;
sine[2173] =63;
sine[2174] =63;
sine[2175] =63;
sine[2176] =63;
sine[2177] =64;
sine[2178] =64;
sine[2179] =64;
sine[2180] =64;
sine[2181] =65;
sine[2182] =65;
sine[2183] =65;
sine[2184] =65;
sine[2185] =66;
sine[2186] =66;
sine[2187] =66;
sine[2188] =66;
sine[2189] =67;
sine[2190] =67;
sine[2191] =67;
sine[2192] =68;
sine[2193] =68;
sine[2194] =68;
sine[2195] =68;
sine[2196] =69;
sine[2197] =69;
sine[2198] =69;
sine[2199] =69;
sine[2200] =70;
sine[2201] =70;
sine[2202] =70;
sine[2203] =70;
sine[2204] =71;
sine[2205] =71;
sine[2206] =71;
sine[2207] =72;
sine[2208] =72;
sine[2209] =72;
sine[2210] =72;
sine[2211] =73;
sine[2212] =73;
sine[2213] =73;
sine[2214] =73;
sine[2215] =74;
sine[2216] =74;
sine[2217] =74;
sine[2218] =75;
sine[2219] =75;
sine[2220] =75;
sine[2221] =75;
sine[2222] =76;
sine[2223] =76;
sine[2224] =76;
sine[2225] =77;
sine[2226] =77;
sine[2227] =77;
sine[2228] =77;
sine[2229] =78;
sine[2230] =78;
sine[2231] =78;
sine[2232] =78;
sine[2233] =79;
sine[2234] =79;
sine[2235] =79;
sine[2236] =80;
sine[2237] =80;
sine[2238] =80;
sine[2239] =80;
sine[2240] =81;
sine[2241] =81;
sine[2242] =81;
sine[2243] =82;
sine[2244] =82;
sine[2245] =82;
sine[2246] =82;
sine[2247] =83;
sine[2248] =83;
sine[2249] =83;
sine[2250] =84;
sine[2251] =84;
sine[2252] =84;
sine[2253] =84;
sine[2254] =85;
sine[2255] =85;
sine[2256] =85;
sine[2257] =86;
sine[2258] =86;
sine[2259] =86;
sine[2260] =87;
sine[2261] =87;
sine[2262] =87;
sine[2263] =87;
sine[2264] =88;
sine[2265] =88;
sine[2266] =88;
sine[2267] =89;
sine[2268] =89;
sine[2269] =89;
sine[2270] =90;
sine[2271] =90;
sine[2272] =90;
sine[2273] =90;
sine[2274] =91;
sine[2275] =91;
sine[2276] =91;
sine[2277] =92;
sine[2278] =92;
sine[2279] =92;
sine[2280] =93;
sine[2281] =93;
sine[2282] =93;
sine[2283] =93;
sine[2284] =94;
sine[2285] =94;
sine[2286] =94;
sine[2287] =95;
sine[2288] =95;
sine[2289] =95;
sine[2290] =96;
sine[2291] =96;
sine[2292] =96;
sine[2293] =96;
sine[2294] =97;
sine[2295] =97;
sine[2296] =97;
sine[2297] =98;
sine[2298] =98;
sine[2299] =98;
sine[2300] =99;
sine[2301] =99;
sine[2302] =99;
sine[2303] =100;
sine[2304] =100;
sine[2305] =100;
sine[2306] =100;
sine[2307] =101;
sine[2308] =101;
sine[2309] =101;
sine[2310] =102;
sine[2311] =102;
sine[2312] =102;
sine[2313] =103;
sine[2314] =103;
sine[2315] =103;
sine[2316] =104;
sine[2317] =104;
sine[2318] =104;
sine[2319] =105;
sine[2320] =105;
sine[2321] =105;
sine[2322] =106;
sine[2323] =106;
sine[2324] =106;
sine[2325] =106;
sine[2326] =107;
sine[2327] =107;
sine[2328] =107;
sine[2329] =108;
sine[2330] =108;
sine[2331] =108;
sine[2332] =109;
sine[2333] =109;
sine[2334] =109;
sine[2335] =110;
sine[2336] =110;
sine[2337] =110;
sine[2338] =111;
sine[2339] =111;
sine[2340] =111;
sine[2341] =112;
sine[2342] =112;
sine[2343] =112;
sine[2344] =113;
sine[2345] =113;
sine[2346] =113;
sine[2347] =114;
sine[2348] =114;
sine[2349] =114;
sine[2350] =115;
sine[2351] =115;
sine[2352] =115;
sine[2353] =116;
sine[2354] =116;
sine[2355] =116;
sine[2356] =116;
sine[2357] =117;
sine[2358] =117;
sine[2359] =117;
sine[2360] =118;
sine[2361] =118;
sine[2362] =118;
sine[2363] =119;
sine[2364] =119;
sine[2365] =119;
sine[2366] =120;
sine[2367] =120;
sine[2368] =120;
sine[2369] =121;
sine[2370] =121;
sine[2371] =121;
sine[2372] =122;
sine[2373] =122;
sine[2374] =122;
sine[2375] =123;
sine[2376] =123;
sine[2377] =123;
sine[2378] =124;
sine[2379] =124;
sine[2380] =124;
sine[2381] =125;
sine[2382] =125;
sine[2383] =125;
sine[2384] =126;
sine[2385] =126;
sine[2386] =127;
sine[2387] =127;
sine[2388] =127;
sine[2389] =128;
sine[2390] =128;
sine[2391] =128;
sine[2392] =129;
sine[2393] =129;
sine[2394] =129;
sine[2395] =130;
sine[2396] =130;
sine[2397] =130;
sine[2398] =131;
sine[2399] =131;
sine[2400] =131;
sine[2401] =132;
sine[2402] =132;
sine[2403] =132;
sine[2404] =133;
sine[2405] =133;
sine[2406] =133;
sine[2407] =134;
sine[2408] =134;
sine[2409] =134;
sine[2410] =135;
sine[2411] =135;
sine[2412] =135;
sine[2413] =136;
sine[2414] =136;
sine[2415] =136;
sine[2416] =137;
sine[2417] =137;
sine[2418] =137;
sine[2419] =138;
sine[2420] =138;
sine[2421] =139;
sine[2422] =139;
sine[2423] =139;
sine[2424] =140;
sine[2425] =140;
sine[2426] =140;
sine[2427] =141;
sine[2428] =141;
sine[2429] =141;
sine[2430] =142;
sine[2431] =142;
sine[2432] =142;
sine[2433] =143;
sine[2434] =143;
sine[2435] =143;
sine[2436] =144;
sine[2437] =144;
sine[2438] =144;
sine[2439] =145;
sine[2440] =145;
sine[2441] =146;
sine[2442] =146;
sine[2443] =146;
sine[2444] =147;
sine[2445] =147;
sine[2446] =147;
sine[2447] =148;
sine[2448] =148;
sine[2449] =148;
sine[2450] =149;
sine[2451] =149;
sine[2452] =149;
sine[2453] =150;
sine[2454] =150;
sine[2455] =151;
sine[2456] =151;
sine[2457] =151;
sine[2458] =152;
sine[2459] =152;
sine[2460] =152;
sine[2461] =153;
sine[2462] =153;
sine[2463] =153;
sine[2464] =154;
sine[2465] =154;
sine[2466] =154;
sine[2467] =155;
sine[2468] =155;
sine[2469] =156;
sine[2470] =156;
sine[2471] =156;
sine[2472] =157;
sine[2473] =157;
sine[2474] =157;
sine[2475] =158;
sine[2476] =158;
sine[2477] =158;
sine[2478] =159;
sine[2479] =159;
sine[2480] =160;
sine[2481] =160;
sine[2482] =160;
sine[2483] =161;
sine[2484] =161;
sine[2485] =161;
sine[2486] =162;
sine[2487] =162;
sine[2488] =162;
sine[2489] =163;
sine[2490] =163;
sine[2491] =164;
sine[2492] =164;
sine[2493] =164;
sine[2494] =165;
sine[2495] =165;
sine[2496] =165;
sine[2497] =166;
sine[2498] =166;
sine[2499] =166;
sine[2500] =167;
sine[2501] =167;
sine[2502] =168;
sine[2503] =168;
sine[2504] =168;
sine[2505] =169;
sine[2506] =169;
sine[2507] =169;
sine[2508] =170;
sine[2509] =170;
sine[2510] =171;
sine[2511] =171;
sine[2512] =171;
sine[2513] =172;
sine[2514] =172;
sine[2515] =172;
sine[2516] =173;
sine[2517] =173;
sine[2518] =173;
sine[2519] =174;
sine[2520] =174;
sine[2521] =175;
sine[2522] =175;
sine[2523] =175;
sine[2524] =176;
sine[2525] =176;
sine[2526] =176;
sine[2527] =177;
sine[2528] =177;
sine[2529] =178;
sine[2530] =178;
sine[2531] =178;
sine[2532] =179;
sine[2533] =179;
sine[2534] =179;
sine[2535] =180;
sine[2536] =180;
sine[2537] =181;
sine[2538] =181;
sine[2539] =181;
sine[2540] =182;
sine[2541] =182;
sine[2542] =182;
sine[2543] =183;
sine[2544] =183;
sine[2545] =184;
sine[2546] =184;
sine[2547] =184;
sine[2548] =185;
sine[2549] =185;
sine[2550] =185;
sine[2551] =186;
sine[2552] =186;
sine[2553] =187;
sine[2554] =187;
sine[2555] =187;
sine[2556] =188;
sine[2557] =188;
sine[2558] =188;
sine[2559] =189;
sine[2560] =189;
sine[2561] =190;
sine[2562] =190;
sine[2563] =190;
sine[2564] =191;
sine[2565] =191;
sine[2566] =192;
sine[2567] =192;
sine[2568] =192;
sine[2569] =193;
sine[2570] =193;
sine[2571] =193;
sine[2572] =194;
sine[2573] =194;
sine[2574] =195;
sine[2575] =195;
sine[2576] =195;
sine[2577] =196;
sine[2578] =196;
sine[2579] =196;
sine[2580] =197;
sine[2581] =197;
sine[2582] =198;
sine[2583] =198;
sine[2584] =198;
sine[2585] =199;
sine[2586] =199;
sine[2587] =200;
sine[2588] =200;
sine[2589] =200;
sine[2590] =201;
sine[2591] =201;
sine[2592] =201;
sine[2593] =202;
sine[2594] =202;
sine[2595] =203;
sine[2596] =203;
sine[2597] =203;
sine[2598] =204;
sine[2599] =204;
sine[2600] =205;
sine[2601] =205;
sine[2602] =205;
sine[2603] =206;
sine[2604] =206;
sine[2605] =206;
sine[2606] =207;
sine[2607] =207;
sine[2608] =208;
sine[2609] =208;
sine[2610] =208;
sine[2611] =209;
sine[2612] =209;
sine[2613] =210;
sine[2614] =210;
sine[2615] =210;
sine[2616] =211;
sine[2617] =211;
sine[2618] =211;
sine[2619] =212;
sine[2620] =212;
sine[2621] =213;
sine[2622] =213;
sine[2623] =213;
sine[2624] =214;
sine[2625] =214;
sine[2626] =215;
sine[2627] =215;
sine[2628] =215;
sine[2629] =216;
sine[2630] =216;
sine[2631] =216;
sine[2632] =217;
sine[2633] =217;
sine[2634] =218;
sine[2635] =218;
sine[2636] =218;
sine[2637] =219;
sine[2638] =219;
sine[2639] =220;
sine[2640] =220;
sine[2641] =220;
sine[2642] =221;
sine[2643] =221;
sine[2644] =222;
sine[2645] =222;
sine[2646] =222;
sine[2647] =223;
sine[2648] =223;
sine[2649] =223;
sine[2650] =224;
sine[2651] =224;
sine[2652] =225;
sine[2653] =225;
sine[2654] =225;
sine[2655] =226;
sine[2656] =226;
sine[2657] =227;
sine[2658] =227;
sine[2659] =227;
sine[2660] =228;
sine[2661] =228;
sine[2662] =229;
sine[2663] =229;
sine[2664] =229;
sine[2665] =230;
sine[2666] =230;
sine[2667] =230;
sine[2668] =231;
sine[2669] =231;
sine[2670] =232;
sine[2671] =232;
sine[2672] =232;
sine[2673] =233;
sine[2674] =233;
sine[2675] =234;
sine[2676] =234;
sine[2677] =234;
sine[2678] =235;
sine[2679] =235;
sine[2680] =236;
sine[2681] =236;
sine[2682] =236;
sine[2683] =237;
sine[2684] =237;
sine[2685] =237;
sine[2686] =238;
sine[2687] =238;
sine[2688] =239;
sine[2689] =239;
sine[2690] =239;
sine[2691] =240;
sine[2692] =240;
sine[2693] =241;
sine[2694] =241;
sine[2695] =241;
sine[2696] =242;
sine[2697] =242;
sine[2698] =243;
sine[2699] =243;
sine[2700] =243;
sine[2701] =244;
sine[2702] =244;
sine[2703] =245;
sine[2704] =245;
sine[2705] =245;
sine[2706] =246;
sine[2707] =246;
sine[2708] =246;
sine[2709] =247;
sine[2710] =247;
sine[2711] =248;
sine[2712] =248;
sine[2713] =248;
sine[2714] =249;
sine[2715] =249;
sine[2716] =250;
sine[2717] =250;
sine[2718] =250;
sine[2719] =251;
sine[2720] =251;
sine[2721] =252;
sine[2722] =252;
sine[2723] =252;
sine[2724] =253;
sine[2725] =253;
sine[2726] =254;
sine[2727] =254;
sine[2728] =254;
sine[2729] =255;
sine[2730] =255;
sine[2731] =256;
sine[2732] =256;
sine[2733] =256;
sine[2734] =257;
sine[2735] =257;
sine[2736] =257;
sine[2737] =258;
sine[2738] =258;
sine[2739] =259;
sine[2740] =259;
sine[2741] =259;
sine[2742] =260;
sine[2743] =260;
sine[2744] =261;
sine[2745] =261;
sine[2746] =261;
sine[2747] =262;
sine[2748] =262;
sine[2749] =263;
sine[2750] =263;
sine[2751] =263;
sine[2752] =264;
sine[2753] =264;
sine[2754] =265;
sine[2755] =265;
sine[2756] =265;
sine[2757] =266;
sine[2758] =266;
sine[2759] =266;
sine[2760] =267;
sine[2761] =267;
sine[2762] =268;
sine[2763] =268;
sine[2764] =268;
sine[2765] =269;
sine[2766] =269;
sine[2767] =270;
sine[2768] =270;
sine[2769] =270;
sine[2770] =271;
sine[2771] =271;
sine[2772] =272;
sine[2773] =272;
sine[2774] =272;
sine[2775] =273;
sine[2776] =273;
sine[2777] =274;
sine[2778] =274;
sine[2779] =274;
sine[2780] =275;
sine[2781] =275;
sine[2782] =275;
sine[2783] =276;
sine[2784] =276;
sine[2785] =277;
sine[2786] =277;
sine[2787] =277;
sine[2788] =278;
sine[2789] =278;
sine[2790] =279;
sine[2791] =279;
sine[2792] =279;
sine[2793] =280;
sine[2794] =280;
sine[2795] =281;
sine[2796] =281;
sine[2797] =281;
sine[2798] =282;
sine[2799] =282;
sine[2800] =282;
sine[2801] =283;
sine[2802] =283;
sine[2803] =284;
sine[2804] =284;
sine[2805] =284;
sine[2806] =285;
sine[2807] =285;
sine[2808] =286;
sine[2809] =286;
sine[2810] =286;
sine[2811] =287;
sine[2812] =287;
sine[2813] =288;
sine[2814] =288;
sine[2815] =288;
sine[2816] =289;
sine[2817] =289;
sine[2818] =289;
sine[2819] =290;
sine[2820] =290;
sine[2821] =291;
sine[2822] =291;
sine[2823] =291;
sine[2824] =292;
sine[2825] =292;
sine[2826] =293;
sine[2827] =293;
sine[2828] =293;
sine[2829] =294;
sine[2830] =294;
sine[2831] =295;
sine[2832] =295;
sine[2833] =295;
sine[2834] =296;
sine[2835] =296;
sine[2836] =296;
sine[2837] =297;
sine[2838] =297;
sine[2839] =298;
sine[2840] =298;
sine[2841] =298;
sine[2842] =299;
sine[2843] =299;
sine[2844] =300;
sine[2845] =300;
sine[2846] =300;
sine[2847] =301;
sine[2848] =301;
sine[2849] =301;
sine[2850] =302;
sine[2851] =302;
sine[2852] =303;
sine[2853] =303;
sine[2854] =303;
sine[2855] =304;
sine[2856] =304;
sine[2857] =305;
sine[2858] =305;
sine[2859] =305;
sine[2860] =306;
sine[2861] =306;
sine[2862] =306;
sine[2863] =307;
sine[2864] =307;
sine[2865] =308;
sine[2866] =308;
sine[2867] =308;
sine[2868] =309;
sine[2869] =309;
sine[2870] =310;
sine[2871] =310;
sine[2872] =310;
sine[2873] =311;
sine[2874] =311;
sine[2875] =311;
sine[2876] =312;
sine[2877] =312;
sine[2878] =313;
sine[2879] =313;
sine[2880] =313;
sine[2881] =314;
sine[2882] =314;
sine[2883] =315;
sine[2884] =315;
sine[2885] =315;
sine[2886] =316;
sine[2887] =316;
sine[2888] =316;
sine[2889] =317;
sine[2890] =317;
sine[2891] =318;
sine[2892] =318;
sine[2893] =318;
sine[2894] =319;
sine[2895] =319;
sine[2896] =319;
sine[2897] =320;
sine[2898] =320;
sine[2899] =321;
sine[2900] =321;
sine[2901] =321;
sine[2902] =322;
sine[2903] =322;
sine[2904] =323;
sine[2905] =323;
sine[2906] =323;
sine[2907] =324;
sine[2908] =324;
sine[2909] =324;
sine[2910] =325;
sine[2911] =325;
sine[2912] =326;
sine[2913] =326;
sine[2914] =326;
sine[2915] =327;
sine[2916] =327;
sine[2917] =327;
sine[2918] =328;
sine[2919] =328;
sine[2920] =329;
sine[2921] =329;
sine[2922] =329;
sine[2923] =330;
sine[2924] =330;
sine[2925] =330;
sine[2926] =331;
sine[2927] =331;
sine[2928] =332;
sine[2929] =332;
sine[2930] =332;
sine[2931] =333;
sine[2932] =333;
sine[2933] =333;
sine[2934] =334;
sine[2935] =334;
sine[2936] =335;
sine[2937] =335;
sine[2938] =335;
sine[2939] =336;
sine[2940] =336;
sine[2941] =336;
sine[2942] =337;
sine[2943] =337;
sine[2944] =338;
sine[2945] =338;
sine[2946] =338;
sine[2947] =339;
sine[2948] =339;
sine[2949] =339;
sine[2950] =340;
sine[2951] =340;
sine[2952] =340;
sine[2953] =341;
sine[2954] =341;
sine[2955] =342;
sine[2956] =342;
sine[2957] =342;
sine[2958] =343;
sine[2959] =343;
sine[2960] =343;
sine[2961] =344;
sine[2962] =344;
sine[2963] =345;
sine[2964] =345;
sine[2965] =345;
sine[2966] =346;
sine[2967] =346;
sine[2968] =346;
sine[2969] =347;
sine[2970] =347;
sine[2971] =347;
sine[2972] =348;
sine[2973] =348;
sine[2974] =349;
sine[2975] =349;
sine[2976] =349;
sine[2977] =350;
sine[2978] =350;
sine[2979] =350;
sine[2980] =351;
sine[2981] =351;
sine[2982] =351;
sine[2983] =352;
sine[2984] =352;
sine[2985] =353;
sine[2986] =353;
sine[2987] =353;
sine[2988] =354;
sine[2989] =354;
sine[2990] =354;
sine[2991] =355;
sine[2992] =355;
sine[2993] =355;
sine[2994] =356;
sine[2995] =356;
sine[2996] =357;
sine[2997] =357;
sine[2998] =357;
sine[2999] =358;
sine[3000] =358;
sine[3001] =358;
sine[3002] =359;
sine[3003] =359;
sine[3004] =359;
sine[3005] =360;
sine[3006] =360;
sine[3007] =360;
sine[3008] =361;
sine[3009] =361;
sine[3010] =362;
sine[3011] =362;
sine[3012] =362;
sine[3013] =363;
sine[3014] =363;
sine[3015] =363;
sine[3016] =364;
sine[3017] =364;
sine[3018] =364;
sine[3019] =365;
sine[3020] =365;
sine[3021] =365;
sine[3022] =366;
sine[3023] =366;
sine[3024] =367;
sine[3025] =367;
sine[3026] =367;
sine[3027] =368;
sine[3028] =368;
sine[3029] =368;
sine[3030] =369;
sine[3031] =369;
sine[3032] =369;
sine[3033] =370;
sine[3034] =370;
sine[3035] =370;
sine[3036] =371;
sine[3037] =371;
sine[3038] =371;
sine[3039] =372;
sine[3040] =372;
sine[3041] =372;
sine[3042] =373;
sine[3043] =373;
sine[3044] =374;
sine[3045] =374;
sine[3046] =374;
sine[3047] =375;
sine[3048] =375;
sine[3049] =375;
sine[3050] =376;
sine[3051] =376;
sine[3052] =376;
sine[3053] =377;
sine[3054] =377;
sine[3055] =377;
sine[3056] =378;
sine[3057] =378;
sine[3058] =378;
sine[3059] =379;
sine[3060] =379;
sine[3061] =379;
sine[3062] =380;
sine[3063] =380;
sine[3064] =380;
sine[3065] =381;
sine[3066] =381;
sine[3067] =381;
sine[3068] =382;
sine[3069] =382;
sine[3070] =382;
sine[3071] =383;
sine[3072] =383;
sine[3073] =383;
sine[3074] =384;
sine[3075] =384;
sine[3076] =384;
sine[3077] =385;
sine[3078] =385;
sine[3079] =386;
sine[3080] =386;
sine[3081] =386;
sine[3082] =387;
sine[3083] =387;
sine[3084] =387;
sine[3085] =388;
sine[3086] =388;
sine[3087] =388;
sine[3088] =389;
sine[3089] =389;
sine[3090] =389;
sine[3091] =390;
sine[3092] =390;
sine[3093] =390;
sine[3094] =391;
sine[3095] =391;
sine[3096] =391;
sine[3097] =392;
sine[3098] =392;
sine[3099] =392;
sine[3100] =393;
sine[3101] =393;
sine[3102] =393;
sine[3103] =394;
sine[3104] =394;
sine[3105] =394;
sine[3106] =395;
sine[3107] =395;
sine[3108] =395;
sine[3109] =395;
sine[3110] =396;
sine[3111] =396;
sine[3112] =396;
sine[3113] =397;
sine[3114] =397;
sine[3115] =397;
sine[3116] =398;
sine[3117] =398;
sine[3118] =398;
sine[3119] =399;
sine[3120] =399;
sine[3121] =399;
sine[3122] =400;
sine[3123] =400;
sine[3124] =400;
sine[3125] =401;
sine[3126] =401;
sine[3127] =401;
sine[3128] =402;
sine[3129] =402;
sine[3130] =402;
sine[3131] =403;
sine[3132] =403;
sine[3133] =403;
sine[3134] =404;
sine[3135] =404;
sine[3136] =404;
sine[3137] =405;
sine[3138] =405;
sine[3139] =405;
sine[3140] =405;
sine[3141] =406;
sine[3142] =406;
sine[3143] =406;
sine[3144] =407;
sine[3145] =407;
sine[3146] =407;
sine[3147] =408;
sine[3148] =408;
sine[3149] =408;
sine[3150] =409;
sine[3151] =409;
sine[3152] =409;
sine[3153] =410;
sine[3154] =410;
sine[3155] =410;
sine[3156] =411;
sine[3157] =411;
sine[3158] =411;
sine[3159] =411;
sine[3160] =412;
sine[3161] =412;
sine[3162] =412;
sine[3163] =413;
sine[3164] =413;
sine[3165] =413;
sine[3166] =414;
sine[3167] =414;
sine[3168] =414;
sine[3169] =415;
sine[3170] =415;
sine[3171] =415;
sine[3172] =415;
sine[3173] =416;
sine[3174] =416;
sine[3175] =416;
sine[3176] =417;
sine[3177] =417;
sine[3178] =417;
sine[3179] =418;
sine[3180] =418;
sine[3181] =418;
sine[3182] =418;
sine[3183] =419;
sine[3184] =419;
sine[3185] =419;
sine[3186] =420;
sine[3187] =420;
sine[3188] =420;
sine[3189] =421;
sine[3190] =421;
sine[3191] =421;
sine[3192] =421;
sine[3193] =422;
sine[3194] =422;
sine[3195] =422;
sine[3196] =423;
sine[3197] =423;
sine[3198] =423;
sine[3199] =424;
sine[3200] =424;
sine[3201] =424;
sine[3202] =424;
sine[3203] =425;
sine[3204] =425;
sine[3205] =425;
sine[3206] =426;
sine[3207] =426;
sine[3208] =426;
sine[3209] =427;
sine[3210] =427;
sine[3211] =427;
sine[3212] =427;
sine[3213] =428;
sine[3214] =428;
sine[3215] =428;
sine[3216] =429;
sine[3217] =429;
sine[3218] =429;
sine[3219] =429;
sine[3220] =430;
sine[3221] =430;
sine[3222] =430;
sine[3223] =431;
sine[3224] =431;
sine[3225] =431;
sine[3226] =431;
sine[3227] =432;
sine[3228] =432;
sine[3229] =432;
sine[3230] =433;
sine[3231] =433;
sine[3232] =433;
sine[3233] =433;
sine[3234] =434;
sine[3235] =434;
sine[3236] =434;
sine[3237] =434;
sine[3238] =435;
sine[3239] =435;
sine[3240] =435;
sine[3241] =436;
sine[3242] =436;
sine[3243] =436;
sine[3244] =436;
sine[3245] =437;
sine[3246] =437;
sine[3247] =437;
sine[3248] =438;
sine[3249] =438;
sine[3250] =438;
sine[3251] =438;
sine[3252] =439;
sine[3253] =439;
sine[3254] =439;
sine[3255] =439;
sine[3256] =440;
sine[3257] =440;
sine[3258] =440;
sine[3259] =441;
sine[3260] =441;
sine[3261] =441;
sine[3262] =441;
sine[3263] =442;
sine[3264] =442;
sine[3265] =442;
sine[3266] =442;
sine[3267] =443;
sine[3268] =443;
sine[3269] =443;
sine[3270] =443;
sine[3271] =444;
sine[3272] =444;
sine[3273] =444;
sine[3274] =445;
sine[3275] =445;
sine[3276] =445;
sine[3277] =445;
sine[3278] =446;
sine[3279] =446;
sine[3280] =446;
sine[3281] =446;
sine[3282] =447;
sine[3283] =447;
sine[3284] =447;
sine[3285] =447;
sine[3286] =448;
sine[3287] =448;
sine[3288] =448;
sine[3289] =448;
sine[3290] =449;
sine[3291] =449;
sine[3292] =449;
sine[3293] =449;
sine[3294] =450;
sine[3295] =450;
sine[3296] =450;
sine[3297] =450;
sine[3298] =451;
sine[3299] =451;
sine[3300] =451;
sine[3301] =452;
sine[3302] =452;
sine[3303] =452;
sine[3304] =452;
sine[3305] =453;
sine[3306] =453;
sine[3307] =453;
sine[3308] =453;
sine[3309] =454;
sine[3310] =454;
sine[3311] =454;
sine[3312] =454;
sine[3313] =454;
sine[3314] =455;
sine[3315] =455;
sine[3316] =455;
sine[3317] =455;
sine[3318] =456;
sine[3319] =456;
sine[3320] =456;
sine[3321] =456;
sine[3322] =457;
sine[3323] =457;
sine[3324] =457;
sine[3325] =457;
sine[3326] =458;
sine[3327] =458;
sine[3328] =458;
sine[3329] =458;
sine[3330] =459;
sine[3331] =459;
sine[3332] =459;
sine[3333] =459;
sine[3334] =460;
sine[3335] =460;
sine[3336] =460;
sine[3337] =460;
sine[3338] =460;
sine[3339] =461;
sine[3340] =461;
sine[3341] =461;
sine[3342] =461;
sine[3343] =462;
sine[3344] =462;
sine[3345] =462;
sine[3346] =462;
sine[3347] =463;
sine[3348] =463;
sine[3349] =463;
sine[3350] =463;
sine[3351] =463;
sine[3352] =464;
sine[3353] =464;
sine[3354] =464;
sine[3355] =464;
sine[3356] =465;
sine[3357] =465;
sine[3358] =465;
sine[3359] =465;
sine[3360] =466;
sine[3361] =466;
sine[3362] =466;
sine[3363] =466;
sine[3364] =466;
sine[3365] =467;
sine[3366] =467;
sine[3367] =467;
sine[3368] =467;
sine[3369] =468;
sine[3370] =468;
sine[3371] =468;
sine[3372] =468;
sine[3373] =468;
sine[3374] =469;
sine[3375] =469;
sine[3376] =469;
sine[3377] =469;
sine[3378] =469;
sine[3379] =470;
sine[3380] =470;
sine[3381] =470;
sine[3382] =470;
sine[3383] =471;
sine[3384] =471;
sine[3385] =471;
sine[3386] =471;
sine[3387] =471;
sine[3388] =472;
sine[3389] =472;
sine[3390] =472;
sine[3391] =472;
sine[3392] =472;
sine[3393] =473;
sine[3394] =473;
sine[3395] =473;
sine[3396] =473;
sine[3397] =473;
sine[3398] =474;
sine[3399] =474;
sine[3400] =474;
sine[3401] =474;
sine[3402] =474;
sine[3403] =475;
sine[3404] =475;
sine[3405] =475;
sine[3406] =475;
sine[3407] =475;
sine[3408] =476;
sine[3409] =476;
sine[3410] =476;
sine[3411] =476;
sine[3412] =476;
sine[3413] =477;
sine[3414] =477;
sine[3415] =477;
sine[3416] =477;
sine[3417] =477;
sine[3418] =478;
sine[3419] =478;
sine[3420] =478;
sine[3421] =478;
sine[3422] =478;
sine[3423] =479;
sine[3424] =479;
sine[3425] =479;
sine[3426] =479;
sine[3427] =479;
sine[3428] =480;
sine[3429] =480;
sine[3430] =480;
sine[3431] =480;
sine[3432] =480;
sine[3433] =480;
sine[3434] =481;
sine[3435] =481;
sine[3436] =481;
sine[3437] =481;
sine[3438] =481;
sine[3439] =482;
sine[3440] =482;
sine[3441] =482;
sine[3442] =482;
sine[3443] =482;
sine[3444] =482;
sine[3445] =483;
sine[3446] =483;
sine[3447] =483;
sine[3448] =483;
sine[3449] =483;
sine[3450] =484;
sine[3451] =484;
sine[3452] =484;
sine[3453] =484;
sine[3454] =484;
sine[3455] =484;
sine[3456] =485;
sine[3457] =485;
sine[3458] =485;
sine[3459] =485;
sine[3460] =485;
sine[3461] =485;
sine[3462] =486;
sine[3463] =486;
sine[3464] =486;
sine[3465] =486;
sine[3466] =486;
sine[3467] =486;
sine[3468] =487;
sine[3469] =487;
sine[3470] =487;
sine[3471] =487;
sine[3472] =487;
sine[3473] =487;
sine[3474] =488;
sine[3475] =488;
sine[3476] =488;
sine[3477] =488;
sine[3478] =488;
sine[3479] =488;
sine[3480] =489;
sine[3481] =489;
sine[3482] =489;
sine[3483] =489;
sine[3484] =489;
sine[3485] =489;
sine[3486] =490;
sine[3487] =490;
sine[3488] =490;
sine[3489] =490;
sine[3490] =490;
sine[3491] =490;
sine[3492] =490;
sine[3493] =491;
sine[3494] =491;
sine[3495] =491;
sine[3496] =491;
sine[3497] =491;
sine[3498] =491;
sine[3499] =492;
sine[3500] =492;
sine[3501] =492;
sine[3502] =492;
sine[3503] =492;
sine[3504] =492;
sine[3505] =492;
sine[3506] =493;
sine[3507] =493;
sine[3508] =493;
sine[3509] =493;
sine[3510] =493;
sine[3511] =493;
sine[3512] =493;
sine[3513] =494;
sine[3514] =494;
sine[3515] =494;
sine[3516] =494;
sine[3517] =494;
sine[3518] =494;
sine[3519] =494;
sine[3520] =495;
sine[3521] =495;
sine[3522] =495;
sine[3523] =495;
sine[3524] =495;
sine[3525] =495;
sine[3526] =495;
sine[3527] =496;
sine[3528] =496;
sine[3529] =496;
sine[3530] =496;
sine[3531] =496;
sine[3532] =496;
sine[3533] =496;
sine[3534] =496;
sine[3535] =497;
sine[3536] =497;
sine[3537] =497;
sine[3538] =497;
sine[3539] =497;
sine[3540] =497;
sine[3541] =497;
sine[3542] =497;
sine[3543] =498;
sine[3544] =498;
sine[3545] =498;
sine[3546] =498;
sine[3547] =498;
sine[3548] =498;
sine[3549] =498;
sine[3550] =498;
sine[3551] =499;
sine[3552] =499;
sine[3553] =499;
sine[3554] =499;
sine[3555] =499;
sine[3556] =499;
sine[3557] =499;
sine[3558] =499;
sine[3559] =500;
sine[3560] =500;
sine[3561] =500;
sine[3562] =500;
sine[3563] =500;
sine[3564] =500;
sine[3565] =500;
sine[3566] =500;
sine[3567] =500;
sine[3568] =501;
sine[3569] =501;
sine[3570] =501;
sine[3571] =501;
sine[3572] =501;
sine[3573] =501;
sine[3574] =501;
sine[3575] =501;
sine[3576] =501;
sine[3577] =502;
sine[3578] =502;
sine[3579] =502;
sine[3580] =502;
sine[3581] =502;
sine[3582] =502;
sine[3583] =502;
sine[3584] =502;
sine[3585] =502;
sine[3586] =502;
sine[3587] =503;
sine[3588] =503;
sine[3589] =503;
sine[3590] =503;
sine[3591] =503;
sine[3592] =503;
sine[3593] =503;
sine[3594] =503;
sine[3595] =503;
sine[3596] =503;
sine[3597] =504;
sine[3598] =504;
sine[3599] =504;
sine[3600] =504;
sine[3601] =504;
sine[3602] =504;
sine[3603] =504;
sine[3604] =504;
sine[3605] =504;
sine[3606] =504;
sine[3607] =504;
sine[3608] =505;
sine[3609] =505;
sine[3610] =505;
sine[3611] =505;
sine[3612] =505;
sine[3613] =505;
sine[3614] =505;
sine[3615] =505;
sine[3616] =505;
sine[3617] =505;
sine[3618] =505;
sine[3619] =505;
sine[3620] =506;
sine[3621] =506;
sine[3622] =506;
sine[3623] =506;
sine[3624] =506;
sine[3625] =506;
sine[3626] =506;
sine[3627] =506;
sine[3628] =506;
sine[3629] =506;
sine[3630] =506;
sine[3631] =506;
sine[3632] =506;
sine[3633] =507;
sine[3634] =507;
sine[3635] =507;
sine[3636] =507;
sine[3637] =507;
sine[3638] =507;
sine[3639] =507;
sine[3640] =507;
sine[3641] =507;
sine[3642] =507;
sine[3643] =507;
sine[3644] =507;
sine[3645] =507;
sine[3646] =507;
sine[3647] =508;
sine[3648] =508;
sine[3649] =508;
sine[3650] =508;
sine[3651] =508;
sine[3652] =508;
sine[3653] =508;
sine[3654] =508;
sine[3655] =508;
sine[3656] =508;
sine[3657] =508;
sine[3658] =508;
sine[3659] =508;
sine[3660] =508;
sine[3661] =508;
sine[3662] =508;
sine[3663] =508;
sine[3664] =509;
sine[3665] =509;
sine[3666] =509;
sine[3667] =509;
sine[3668] =509;
sine[3669] =509;
sine[3670] =509;
sine[3671] =509;
sine[3672] =509;
sine[3673] =509;
sine[3674] =509;
sine[3675] =509;
sine[3676] =509;
sine[3677] =509;
sine[3678] =509;
sine[3679] =509;
sine[3680] =509;
sine[3681] =509;
sine[3682] =509;
sine[3683] =509;
sine[3684] =509;
sine[3685] =510;
sine[3686] =510;
sine[3687] =510;
sine[3688] =510;
sine[3689] =510;
sine[3690] =510;
sine[3691] =510;
sine[3692] =510;
sine[3693] =510;
sine[3694] =510;
sine[3695] =510;
sine[3696] =510;
sine[3697] =510;
sine[3698] =510;
sine[3699] =510;
sine[3700] =510;
sine[3701] =510;
sine[3702] =510;
sine[3703] =510;
sine[3704] =510;
sine[3705] =510;
sine[3706] =510;
sine[3707] =510;
sine[3708] =510;
sine[3709] =510;
sine[3710] =510;
sine[3711] =510;
sine[3712] =510;
sine[3713] =510;
sine[3714] =510;
sine[3715] =511;
sine[3716] =511;
sine[3717] =511;
sine[3718] =511;
sine[3719] =511;
sine[3720] =511;
sine[3721] =511;
sine[3722] =511;
sine[3723] =511;
sine[3724] =511;
sine[3725] =511;
sine[3726] =511;
sine[3727] =511;
sine[3728] =511;
sine[3729] =511;
sine[3730] =511;
sine[3731] =511;
sine[3732] =511;
sine[3733] =511;
sine[3734] =511;
sine[3735] =511;
sine[3736] =511;
sine[3737] =511;
sine[3738] =511;
sine[3739] =511;
sine[3740] =511;
sine[3741] =511;
sine[3742] =511;
sine[3743] =511;
sine[3744] =511;
sine[3745] =511;
sine[3746] =511;
sine[3747] =511;
sine[3748] =511;
sine[3749] =511;
sine[3750] =511;
sine[3751] =511;
sine[3752] =511;
sine[3753] =511;
sine[3754] =511;
sine[3755] =511;
sine[3756] =511;
sine[3757] =511;
sine[3758] =511;
sine[3759] =511;
sine[3760] =511;
sine[3761] =511;
sine[3762] =511;
sine[3763] =511;
sine[3764] =511;
sine[3765] =511;
sine[3766] =511;
sine[3767] =511;
sine[3768] =511;
sine[3769] =511;
sine[3770] =511;
sine[3771] =511;
sine[3772] =511;
sine[3773] =511;
sine[3774] =511;
sine[3775] =511;
sine[3776] =511;
sine[3777] =511;
sine[3778] =511;
sine[3779] =511;
sine[3780] =511;
sine[3781] =511;
sine[3782] =511;
sine[3783] =511;
sine[3784] =511;
sine[3785] =511;
sine[3786] =511;
sine[3787] =511;
sine[3788] =511;
sine[3789] =511;
sine[3790] =511;
sine[3791] =511;
sine[3792] =511;
sine[3793] =511;
sine[3794] =511;
sine[3795] =511;
sine[3796] =510;
sine[3797] =510;
sine[3798] =510;
sine[3799] =510;
sine[3800] =510;
sine[3801] =510;
sine[3802] =510;
sine[3803] =510;
sine[3804] =510;
sine[3805] =510;
sine[3806] =510;
sine[3807] =510;
sine[3808] =510;
sine[3809] =510;
sine[3810] =510;
sine[3811] =510;
sine[3812] =510;
sine[3813] =510;
sine[3814] =510;
sine[3815] =510;
sine[3816] =510;
sine[3817] =510;
sine[3818] =510;
sine[3819] =510;
sine[3820] =510;
sine[3821] =510;
sine[3822] =510;
sine[3823] =510;
sine[3824] =510;
sine[3825] =510;
sine[3826] =509;
sine[3827] =509;
sine[3828] =509;
sine[3829] =509;
sine[3830] =509;
sine[3831] =509;
sine[3832] =509;
sine[3833] =509;
sine[3834] =509;
sine[3835] =509;
sine[3836] =509;
sine[3837] =509;
sine[3838] =509;
sine[3839] =509;
sine[3840] =509;
sine[3841] =509;
sine[3842] =509;
sine[3843] =509;
sine[3844] =509;
sine[3845] =509;
sine[3846] =509;
sine[3847] =508;
sine[3848] =508;
sine[3849] =508;
sine[3850] =508;
sine[3851] =508;
sine[3852] =508;
sine[3853] =508;
sine[3854] =508;
sine[3855] =508;
sine[3856] =508;
sine[3857] =508;
sine[3858] =508;
sine[3859] =508;
sine[3860] =508;
sine[3861] =508;
sine[3862] =508;
sine[3863] =508;
sine[3864] =507;
sine[3865] =507;
sine[3866] =507;
sine[3867] =507;
sine[3868] =507;
sine[3869] =507;
sine[3870] =507;
sine[3871] =507;
sine[3872] =507;
sine[3873] =507;
sine[3874] =507;
sine[3875] =507;
sine[3876] =507;
sine[3877] =507;
sine[3878] =506;
sine[3879] =506;
sine[3880] =506;
sine[3881] =506;
sine[3882] =506;
sine[3883] =506;
sine[3884] =506;
sine[3885] =506;
sine[3886] =506;
sine[3887] =506;
sine[3888] =506;
sine[3889] =506;
sine[3890] =506;
sine[3891] =505;
sine[3892] =505;
sine[3893] =505;
sine[3894] =505;
sine[3895] =505;
sine[3896] =505;
sine[3897] =505;
sine[3898] =505;
sine[3899] =505;
sine[3900] =505;
sine[3901] =505;
sine[3902] =505;
sine[3903] =504;
sine[3904] =504;
sine[3905] =504;
sine[3906] =504;
sine[3907] =504;
sine[3908] =504;
sine[3909] =504;
sine[3910] =504;
sine[3911] =504;
sine[3912] =504;
sine[3913] =504;
sine[3914] =503;
sine[3915] =503;
sine[3916] =503;
sine[3917] =503;
sine[3918] =503;
sine[3919] =503;
sine[3920] =503;
sine[3921] =503;
sine[3922] =503;
sine[3923] =503;
sine[3924] =502;
sine[3925] =502;
sine[3926] =502;
sine[3927] =502;
sine[3928] =502;
sine[3929] =502;
sine[3930] =502;
sine[3931] =502;
sine[3932] =502;
sine[3933] =502;
sine[3934] =501;
sine[3935] =501;
sine[3936] =501;
sine[3937] =501;
sine[3938] =501;
sine[3939] =501;
sine[3940] =501;
sine[3941] =501;
sine[3942] =501;
sine[3943] =500;
sine[3944] =500;
sine[3945] =500;
sine[3946] =500;
sine[3947] =500;
sine[3948] =500;
sine[3949] =500;
sine[3950] =500;
sine[3951] =500;
sine[3952] =499;
sine[3953] =499;
sine[3954] =499;
sine[3955] =499;
sine[3956] =499;
sine[3957] =499;
sine[3958] =499;
sine[3959] =499;
sine[3960] =498;
sine[3961] =498;
sine[3962] =498;
sine[3963] =498;
sine[3964] =498;
sine[3965] =498;
sine[3966] =498;
sine[3967] =498;
sine[3968] =497;
sine[3969] =497;
sine[3970] =497;
sine[3971] =497;
sine[3972] =497;
sine[3973] =497;
sine[3974] =497;
sine[3975] =497;
sine[3976] =496;
sine[3977] =496;
sine[3978] =496;
sine[3979] =496;
sine[3980] =496;
sine[3981] =496;
sine[3982] =496;
sine[3983] =496;
sine[3984] =495;
sine[3985] =495;
sine[3986] =495;
sine[3987] =495;
sine[3988] =495;
sine[3989] =495;
sine[3990] =495;
sine[3991] =494;
sine[3992] =494;
sine[3993] =494;
sine[3994] =494;
sine[3995] =494;
sine[3996] =494;
sine[3997] =494;
sine[3998] =493;
sine[3999] =493;
sine[4000] =493;
sine[4001] =493;
sine[4002] =493;
sine[4003] =493;
sine[4004] =493;
sine[4005] =492;
sine[4006] =492;
sine[4007] =492;
sine[4008] =492;
sine[4009] =492;
sine[4010] =492;
sine[4011] =492;
sine[4012] =491;
sine[4013] =491;
sine[4014] =491;
sine[4015] =491;
sine[4016] =491;
sine[4017] =491;
sine[4018] =490;
sine[4019] =490;
sine[4020] =490;
sine[4021] =490;
sine[4022] =490;
sine[4023] =490;
sine[4024] =490;
sine[4025] =489;
sine[4026] =489;
sine[4027] =489;
sine[4028] =489;
sine[4029] =489;
sine[4030] =489;
sine[4031] =488;
sine[4032] =488;
sine[4033] =488;
sine[4034] =488;
sine[4035] =488;
sine[4036] =488;
sine[4037] =487;
sine[4038] =487;
sine[4039] =487;
sine[4040] =487;
sine[4041] =487;
sine[4042] =487;
sine[4043] =486;
sine[4044] =486;
sine[4045] =486;
sine[4046] =486;
sine[4047] =486;
sine[4048] =486;
sine[4049] =485;
sine[4050] =485;
sine[4051] =485;
sine[4052] =485;
sine[4053] =485;
sine[4054] =485;
sine[4055] =484;
sine[4056] =484;
sine[4057] =484;
sine[4058] =484;
sine[4059] =484;
sine[4060] =484;
sine[4061] =483;
sine[4062] =483;
sine[4063] =483;
sine[4064] =483;
sine[4065] =483;
sine[4066] =482;
sine[4067] =482;
sine[4068] =482;
sine[4069] =482;
sine[4070] =482;
sine[4071] =482;
sine[4072] =481;
sine[4073] =481;
sine[4074] =481;
sine[4075] =481;
sine[4076] =481;
sine[4077] =480;
sine[4078] =480;
sine[4079] =480;
sine[4080] =480;
sine[4081] =480;
sine[4082] =480;
sine[4083] =479;
sine[4084] =479;
sine[4085] =479;
sine[4086] =479;
sine[4087] =479;
sine[4088] =478;
sine[4089] =478;
sine[4090] =478;
sine[4091] =478;
sine[4092] =478;
sine[4093] =477;
sine[4094] =477;
sine[4095] =477;
    end
        always@ (posedge(Clk))
    begin
        data_out_2 = sine[j];
        j = j+ 1;
        if(j == 4095)
            j = 0;
    end
endmodule