module LUT_method_1(Clk,reset,data_out_1);
       input Clk,reset;
       output reg [11:0] data_out_1;
       reg [20:0] counter; 
       reg [11:0] sine [0:4095];
       integer i;  
     initial begin
        i = 0;

sine[0] =256;
sine[1] =256;
sine[2] =256;
sine[3] =257;
sine[4] =257;
sine[5] =257;
sine[6] =258;
sine[7] =258;
sine[8] =259;
sine[9] =259;
sine[10] =259;
sine[11] =260;
sine[12] =260;
sine[13] =261;
sine[14] =261;
sine[15] =261;
sine[16] =262;
sine[17] =262;
sine[18] =263;
sine[19] =263;
sine[20] =263;
sine[21] =264;
sine[22] =264;
sine[23] =265;
sine[24] =265;
sine[25] =265;
sine[26] =266;
sine[27] =266;
sine[28] =266;
sine[29] =267;
sine[30] =267;
sine[31] =268;
sine[32] =268;
sine[33] =268;
sine[34] =269;
sine[35] =269;
sine[36] =270;
sine[37] =270;
sine[38] =270;
sine[39] =271;
sine[40] =271;
sine[41] =272;
sine[42] =272;
sine[43] =272;
sine[44] =273;
sine[45] =273;
sine[46] =274;
sine[47] =274;
sine[48] =274;
sine[49] =275;
sine[50] =275;
sine[51] =275;
sine[52] =276;
sine[53] =276;
sine[54] =277;
sine[55] =277;
sine[56] =277;
sine[57] =278;
sine[58] =278;
sine[59] =279;
sine[60] =279;
sine[61] =279;
sine[62] =280;
sine[63] =280;
sine[64] =281;
sine[65] =281;
sine[66] =281;
sine[67] =282;
sine[68] =282;
sine[69] =282;
sine[70] =283;
sine[71] =283;
sine[72] =284;
sine[73] =284;
sine[74] =284;
sine[75] =285;
sine[76] =285;
sine[77] =286;
sine[78] =286;
sine[79] =286;
sine[80] =287;
sine[81] =287;
sine[82] =288;
sine[83] =288;
sine[84] =288;
sine[85] =289;
sine[86] =289;
sine[87] =289;
sine[88] =290;
sine[89] =290;
sine[90] =291;
sine[91] =291;
sine[92] =291;
sine[93] =292;
sine[94] =292;
sine[95] =293;
sine[96] =293;
sine[97] =293;
sine[98] =294;
sine[99] =294;
sine[100] =295;
sine[101] =295;
sine[102] =295;
sine[103] =296;
sine[104] =296;
sine[105] =296;
sine[106] =297;
sine[107] =297;
sine[108] =298;
sine[109] =298;
sine[110] =298;
sine[111] =299;
sine[112] =299;
sine[113] =300;
sine[114] =300;
sine[115] =300;
sine[116] =301;
sine[117] =301;
sine[118] =301;
sine[119] =302;
sine[120] =302;
sine[121] =303;
sine[122] =303;
sine[123] =303;
sine[124] =304;
sine[125] =304;
sine[126] =305;
sine[127] =305;
sine[128] =305;
sine[129] =306;
sine[130] =306;
sine[131] =306;
sine[132] =307;
sine[133] =307;
sine[134] =308;
sine[135] =308;
sine[136] =308;
sine[137] =309;
sine[138] =309;
sine[139] =310;
sine[140] =310;
sine[141] =310;
sine[142] =311;
sine[143] =311;
sine[144] =311;
sine[145] =312;
sine[146] =312;
sine[147] =313;
sine[148] =313;
sine[149] =313;
sine[150] =314;
sine[151] =314;
sine[152] =315;
sine[153] =315;
sine[154] =315;
sine[155] =316;
sine[156] =316;
sine[157] =316;
sine[158] =317;
sine[159] =317;
sine[160] =318;
sine[161] =318;
sine[162] =318;
sine[163] =319;
sine[164] =319;
sine[165] =319;
sine[166] =320;
sine[167] =320;
sine[168] =321;
sine[169] =321;
sine[170] =321;
sine[171] =322;
sine[172] =322;
sine[173] =323;
sine[174] =323;
sine[175] =323;
sine[176] =324;
sine[177] =324;
sine[178] =324;
sine[179] =325;
sine[180] =325;
sine[181] =326;
sine[182] =326;
sine[183] =326;
sine[184] =327;
sine[185] =327;
sine[186] =327;
sine[187] =328;
sine[188] =328;
sine[189] =329;
sine[190] =329;
sine[191] =329;
sine[192] =330;
sine[193] =330;
sine[194] =330;
sine[195] =331;
sine[196] =331;
sine[197] =332;
sine[198] =332;
sine[199] =332;
sine[200] =333;
sine[201] =333;
sine[202] =333;
sine[203] =334;
sine[204] =334;
sine[205] =335;
sine[206] =335;
sine[207] =335;
sine[208] =336;
sine[209] =336;
sine[210] =336;
sine[211] =337;
sine[212] =337;
sine[213] =338;
sine[214] =338;
sine[215] =338;
sine[216] =339;
sine[217] =339;
sine[218] =339;
sine[219] =340;
sine[220] =340;
sine[221] =340;
sine[222] =341;
sine[223] =341;
sine[224] =342;
sine[225] =342;
sine[226] =342;
sine[227] =343;
sine[228] =343;
sine[229] =343;
sine[230] =344;
sine[231] =344;
sine[232] =345;
sine[233] =345;
sine[234] =345;
sine[235] =346;
sine[236] =346;
sine[237] =346;
sine[238] =347;
sine[239] =347;
sine[240] =347;
sine[241] =348;
sine[242] =348;
sine[243] =349;
sine[244] =349;
sine[245] =349;
sine[246] =350;
sine[247] =350;
sine[248] =350;
sine[249] =351;
sine[250] =351;
sine[251] =351;
sine[252] =352;
sine[253] =352;
sine[254] =353;
sine[255] =353;
sine[256] =353;
sine[257] =354;
sine[258] =354;
sine[259] =354;
sine[260] =355;
sine[261] =355;
sine[262] =355;
sine[263] =356;
sine[264] =356;
sine[265] =357;
sine[266] =357;
sine[267] =357;
sine[268] =358;
sine[269] =358;
sine[270] =358;
sine[271] =359;
sine[272] =359;
sine[273] =359;
sine[274] =360;
sine[275] =360;
sine[276] =360;
sine[277] =361;
sine[278] =361;
sine[279] =362;
sine[280] =362;
sine[281] =362;
sine[282] =363;
sine[283] =363;
sine[284] =363;
sine[285] =364;
sine[286] =364;
sine[287] =364;
sine[288] =365;
sine[289] =365;
sine[290] =365;
sine[291] =366;
sine[292] =366;
sine[293] =367;
sine[294] =367;
sine[295] =367;
sine[296] =368;
sine[297] =368;
sine[298] =368;
sine[299] =369;
sine[300] =369;
sine[301] =369;
sine[302] =370;
sine[303] =370;
sine[304] =370;
sine[305] =371;
sine[306] =371;
sine[307] =371;
sine[308] =372;
sine[309] =372;
sine[310] =372;
sine[311] =373;
sine[312] =373;
sine[313] =374;
sine[314] =374;
sine[315] =374;
sine[316] =375;
sine[317] =375;
sine[318] =375;
sine[319] =376;
sine[320] =376;
sine[321] =376;
sine[322] =377;
sine[323] =377;
sine[324] =377;
sine[325] =378;
sine[326] =378;
sine[327] =378;
sine[328] =379;
sine[329] =379;
sine[330] =379;
sine[331] =380;
sine[332] =380;
sine[333] =380;
sine[334] =381;
sine[335] =381;
sine[336] =381;
sine[337] =382;
sine[338] =382;
sine[339] =382;
sine[340] =383;
sine[341] =383;
sine[342] =383;
sine[343] =384;
sine[344] =384;
sine[345] =384;
sine[346] =385;
sine[347] =385;
sine[348] =386;
sine[349] =386;
sine[350] =386;
sine[351] =387;
sine[352] =387;
sine[353] =387;
sine[354] =388;
sine[355] =388;
sine[356] =388;
sine[357] =389;
sine[358] =389;
sine[359] =389;
sine[360] =390;
sine[361] =390;
sine[362] =390;
sine[363] =391;
sine[364] =391;
sine[365] =391;
sine[366] =392;
sine[367] =392;
sine[368] =392;
sine[369] =393;
sine[370] =393;
sine[371] =393;
sine[372] =394;
sine[373] =394;
sine[374] =394;
sine[375] =395;
sine[376] =395;
sine[377] =395;
sine[378] =395;
sine[379] =396;
sine[380] =396;
sine[381] =396;
sine[382] =397;
sine[383] =397;
sine[384] =397;
sine[385] =398;
sine[386] =398;
sine[387] =398;
sine[388] =399;
sine[389] =399;
sine[390] =399;
sine[391] =400;
sine[392] =400;
sine[393] =400;
sine[394] =401;
sine[395] =401;
sine[396] =401;
sine[397] =402;
sine[398] =402;
sine[399] =402;
sine[400] =403;
sine[401] =403;
sine[402] =403;
sine[403] =404;
sine[404] =404;
sine[405] =404;
sine[406] =405;
sine[407] =405;
sine[408] =405;
sine[409] =405;
sine[410] =406;
sine[411] =406;
sine[412] =406;
sine[413] =407;
sine[414] =407;
sine[415] =407;
sine[416] =408;
sine[417] =408;
sine[418] =408;
sine[419] =409;
sine[420] =409;
sine[421] =409;
sine[422] =410;
sine[423] =410;
sine[424] =410;
sine[425] =411;
sine[426] =411;
sine[427] =411;
sine[428] =411;
sine[429] =412;
sine[430] =412;
sine[431] =412;
sine[432] =413;
sine[433] =413;
sine[434] =413;
sine[435] =414;
sine[436] =414;
sine[437] =414;
sine[438] =415;
sine[439] =415;
sine[440] =415;
sine[441] =415;
sine[442] =416;
sine[443] =416;
sine[444] =416;
sine[445] =417;
sine[446] =417;
sine[447] =417;
sine[448] =418;
sine[449] =418;
sine[450] =418;
sine[451] =418;
sine[452] =419;
sine[453] =419;
sine[454] =419;
sine[455] =420;
sine[456] =420;
sine[457] =420;
sine[458] =421;
sine[459] =421;
sine[460] =421;
sine[461] =421;
sine[462] =422;
sine[463] =422;
sine[464] =422;
sine[465] =423;
sine[466] =423;
sine[467] =423;
sine[468] =424;
sine[469] =424;
sine[470] =424;
sine[471] =424;
sine[472] =425;
sine[473] =425;
sine[474] =425;
sine[475] =426;
sine[476] =426;
sine[477] =426;
sine[478] =427;
sine[479] =427;
sine[480] =427;
sine[481] =427;
sine[482] =428;
sine[483] =428;
sine[484] =428;
sine[485] =429;
sine[486] =429;
sine[487] =429;
sine[488] =429;
sine[489] =430;
sine[490] =430;
sine[491] =430;
sine[492] =431;
sine[493] =431;
sine[494] =431;
sine[495] =431;
sine[496] =432;
sine[497] =432;
sine[498] =432;
sine[499] =433;
sine[500] =433;
sine[501] =433;
sine[502] =433;
sine[503] =434;
sine[504] =434;
sine[505] =434;
sine[506] =434;
sine[507] =435;
sine[508] =435;
sine[509] =435;
sine[510] =436;
sine[511] =436;
sine[512] =436;
sine[513] =436;
sine[514] =437;
sine[515] =437;
sine[516] =437;
sine[517] =438;
sine[518] =438;
sine[519] =438;
sine[520] =438;
sine[521] =439;
sine[522] =439;
sine[523] =439;
sine[524] =439;
sine[525] =440;
sine[526] =440;
sine[527] =440;
sine[528] =441;
sine[529] =441;
sine[530] =441;
sine[531] =441;
sine[532] =442;
sine[533] =442;
sine[534] =442;
sine[535] =442;
sine[536] =443;
sine[537] =443;
sine[538] =443;
sine[539] =443;
sine[540] =444;
sine[541] =444;
sine[542] =444;
sine[543] =445;
sine[544] =445;
sine[545] =445;
sine[546] =445;
sine[547] =446;
sine[548] =446;
sine[549] =446;
sine[550] =446;
sine[551] =447;
sine[552] =447;
sine[553] =447;
sine[554] =447;
sine[555] =448;
sine[556] =448;
sine[557] =448;
sine[558] =448;
sine[559] =449;
sine[560] =449;
sine[561] =449;
sine[562] =449;
sine[563] =450;
sine[564] =450;
sine[565] =450;
sine[566] =450;
sine[567] =451;
sine[568] =451;
sine[569] =451;
sine[570] =452;
sine[571] =452;
sine[572] =452;
sine[573] =452;
sine[574] =453;
sine[575] =453;
sine[576] =453;
sine[577] =453;
sine[578] =454;
sine[579] =454;
sine[580] =454;
sine[581] =454;
sine[582] =454;
sine[583] =455;
sine[584] =455;
sine[585] =455;
sine[586] =455;
sine[587] =456;
sine[588] =456;
sine[589] =456;
sine[590] =456;
sine[591] =457;
sine[592] =457;
sine[593] =457;
sine[594] =457;
sine[595] =458;
sine[596] =458;
sine[597] =458;
sine[598] =458;
sine[599] =459;
sine[600] =459;
sine[601] =459;
sine[602] =459;
sine[603] =460;
sine[604] =460;
sine[605] =460;
sine[606] =460;
sine[607] =460;
sine[608] =461;
sine[609] =461;
sine[610] =461;
sine[611] =461;
sine[612] =462;
sine[613] =462;
sine[614] =462;
sine[615] =462;
sine[616] =463;
sine[617] =463;
sine[618] =463;
sine[619] =463;
sine[620] =463;
sine[621] =464;
sine[622] =464;
sine[623] =464;
sine[624] =464;
sine[625] =465;
sine[626] =465;
sine[627] =465;
sine[628] =465;
sine[629] =466;
sine[630] =466;
sine[631] =466;
sine[632] =466;
sine[633] =466;
sine[634] =467;
sine[635] =467;
sine[636] =467;
sine[637] =467;
sine[638] =468;
sine[639] =468;
sine[640] =468;
sine[641] =468;
sine[642] =468;
sine[643] =469;
sine[644] =469;
sine[645] =469;
sine[646] =469;
sine[647] =469;
sine[648] =470;
sine[649] =470;
sine[650] =470;
sine[651] =470;
sine[652] =471;
sine[653] =471;
sine[654] =471;
sine[655] =471;
sine[656] =471;
sine[657] =472;
sine[658] =472;
sine[659] =472;
sine[660] =472;
sine[661] =472;
sine[662] =473;
sine[663] =473;
sine[664] =473;
sine[665] =473;
sine[666] =473;
sine[667] =474;
sine[668] =474;
sine[669] =474;
sine[670] =474;
sine[671] =474;
sine[672] =475;
sine[673] =475;
sine[674] =475;
sine[675] =475;
sine[676] =475;
sine[677] =476;
sine[678] =476;
sine[679] =476;
sine[680] =476;
sine[681] =476;
sine[682] =477;
sine[683] =477;
sine[684] =477;
sine[685] =477;
sine[686] =477;
sine[687] =478;
sine[688] =478;
sine[689] =478;
sine[690] =478;
sine[691] =478;
sine[692] =479;
sine[693] =479;
sine[694] =479;
sine[695] =479;
sine[696] =479;
sine[697] =480;
sine[698] =480;
sine[699] =480;
sine[700] =480;
sine[701] =480;
sine[702] =480;
sine[703] =481;
sine[704] =481;
sine[705] =481;
sine[706] =481;
sine[707] =481;
sine[708] =482;
sine[709] =482;
sine[710] =482;
sine[711] =482;
sine[712] =482;
sine[713] =482;
sine[714] =483;
sine[715] =483;
sine[716] =483;
sine[717] =483;
sine[718] =483;
sine[719] =484;
sine[720] =484;
sine[721] =484;
sine[722] =484;
sine[723] =484;
sine[724] =484;
sine[725] =485;
sine[726] =485;
sine[727] =485;
sine[728] =485;
sine[729] =485;
sine[730] =485;
sine[731] =486;
sine[732] =486;
sine[733] =486;
sine[734] =486;
sine[735] =486;
sine[736] =486;
sine[737] =487;
sine[738] =487;
sine[739] =487;
sine[740] =487;
sine[741] =487;
sine[742] =487;
sine[743] =488;
sine[744] =488;
sine[745] =488;
sine[746] =488;
sine[747] =488;
sine[748] =488;
sine[749] =489;
sine[750] =489;
sine[751] =489;
sine[752] =489;
sine[753] =489;
sine[754] =489;
sine[755] =490;
sine[756] =490;
sine[757] =490;
sine[758] =490;
sine[759] =490;
sine[760] =490;
sine[761] =490;
sine[762] =491;
sine[763] =491;
sine[764] =491;
sine[765] =491;
sine[766] =491;
sine[767] =491;
sine[768] =492;
sine[769] =492;
sine[770] =492;
sine[771] =492;
sine[772] =492;
sine[773] =492;
sine[774] =492;
sine[775] =493;
sine[776] =493;
sine[777] =493;
sine[778] =493;
sine[779] =493;
sine[780] =493;
sine[781] =493;
sine[782] =494;
sine[783] =494;
sine[784] =494;
sine[785] =494;
sine[786] =494;
sine[787] =494;
sine[788] =494;
sine[789] =495;
sine[790] =495;
sine[791] =495;
sine[792] =495;
sine[793] =495;
sine[794] =495;
sine[795] =495;
sine[796] =496;
sine[797] =496;
sine[798] =496;
sine[799] =496;
sine[800] =496;
sine[801] =496;
sine[802] =496;
sine[803] =496;
sine[804] =497;
sine[805] =497;
sine[806] =497;
sine[807] =497;
sine[808] =497;
sine[809] =497;
sine[810] =497;
sine[811] =497;
sine[812] =498;
sine[813] =498;
sine[814] =498;
sine[815] =498;
sine[816] =498;
sine[817] =498;
sine[818] =498;
sine[819] =498;
sine[820] =499;
sine[821] =499;
sine[822] =499;
sine[823] =499;
sine[824] =499;
sine[825] =499;
sine[826] =499;
sine[827] =499;
sine[828] =500;
sine[829] =500;
sine[830] =500;
sine[831] =500;
sine[832] =500;
sine[833] =500;
sine[834] =500;
sine[835] =500;
sine[836] =500;
sine[837] =501;
sine[838] =501;
sine[839] =501;
sine[840] =501;
sine[841] =501;
sine[842] =501;
sine[843] =501;
sine[844] =501;
sine[845] =501;
sine[846] =502;
sine[847] =502;
sine[848] =502;
sine[849] =502;
sine[850] =502;
sine[851] =502;
sine[852] =502;
sine[853] =502;
sine[854] =502;
sine[855] =502;
sine[856] =503;
sine[857] =503;
sine[858] =503;
sine[859] =503;
sine[860] =503;
sine[861] =503;
sine[862] =503;
sine[863] =503;
sine[864] =503;
sine[865] =503;
sine[866] =504;
sine[867] =504;
sine[868] =504;
sine[869] =504;
sine[870] =504;
sine[871] =504;
sine[872] =504;
sine[873] =504;
sine[874] =504;
sine[875] =504;
sine[876] =504;
sine[877] =505;
sine[878] =505;
sine[879] =505;
sine[880] =505;
sine[881] =505;
sine[882] =505;
sine[883] =505;
sine[884] =505;
sine[885] =505;
sine[886] =505;
sine[887] =505;
sine[888] =505;
sine[889] =506;
sine[890] =506;
sine[891] =506;
sine[892] =506;
sine[893] =506;
sine[894] =506;
sine[895] =506;
sine[896] =506;
sine[897] =506;
sine[898] =506;
sine[899] =506;
sine[900] =506;
sine[901] =506;
sine[902] =507;
sine[903] =507;
sine[904] =507;
sine[905] =507;
sine[906] =507;
sine[907] =507;
sine[908] =507;
sine[909] =507;
sine[910] =507;
sine[911] =507;
sine[912] =507;
sine[913] =507;
sine[914] =507;
sine[915] =507;
sine[916] =508;
sine[917] =508;
sine[918] =508;
sine[919] =508;
sine[920] =508;
sine[921] =508;
sine[922] =508;
sine[923] =508;
sine[924] =508;
sine[925] =508;
sine[926] =508;
sine[927] =508;
sine[928] =508;
sine[929] =508;
sine[930] =508;
sine[931] =508;
sine[932] =508;
sine[933] =509;
sine[934] =509;
sine[935] =509;
sine[936] =509;
sine[937] =509;
sine[938] =509;
sine[939] =509;
sine[940] =509;
sine[941] =509;
sine[942] =509;
sine[943] =509;
sine[944] =509;
sine[945] =509;
sine[946] =509;
sine[947] =509;
sine[948] =509;
sine[949] =509;
sine[950] =509;
sine[951] =509;
sine[952] =509;
sine[953] =509;
sine[954] =510;
sine[955] =510;
sine[956] =510;
sine[957] =510;
sine[958] =510;
sine[959] =510;
sine[960] =510;
sine[961] =510;
sine[962] =510;
sine[963] =510;
sine[964] =510;
sine[965] =510;
sine[966] =510;
sine[967] =510;
sine[968] =510;
sine[969] =510;
sine[970] =510;
sine[971] =510;
sine[972] =510;
sine[973] =510;
sine[974] =510;
sine[975] =510;
sine[976] =510;
sine[977] =510;
sine[978] =510;
sine[979] =510;
sine[980] =510;
sine[981] =510;
sine[982] =510;
sine[983] =510;
sine[984] =511;
sine[985] =511;
sine[986] =511;
sine[987] =511;
sine[988] =511;
sine[989] =511;
sine[990] =511;
sine[991] =511;
sine[992] =511;
sine[993] =511;
sine[994] =511;
sine[995] =511;
sine[996] =511;
sine[997] =511;
sine[998] =511;
sine[999] =511;
sine[1000] =511;
sine[1001] =511;
sine[1002] =511;
sine[1003] =511;
sine[1004] =511;
sine[1005] =511;
sine[1006] =511;
sine[1007] =511;
sine[1008] =511;
sine[1009] =511;
sine[1010] =511;
sine[1011] =511;
sine[1012] =511;
sine[1013] =511;
sine[1014] =511;
sine[1015] =511;
sine[1016] =511;
sine[1017] =511;
sine[1018] =511;
sine[1019] =511;
sine[1020] =511;
sine[1021] =511;
sine[1022] =511;
sine[1023] =511;
sine[1024] =511;
sine[1025] =511;
sine[1026] =511;
sine[1027] =511;
sine[1028] =511;
sine[1029] =511;
sine[1030] =511;
sine[1031] =511;
sine[1032] =511;
sine[1033] =511;
sine[1034] =511;
sine[1035] =511;
sine[1036] =511;
sine[1037] =511;
sine[1038] =511;
sine[1039] =511;
sine[1040] =511;
sine[1041] =511;
sine[1042] =511;
sine[1043] =511;
sine[1044] =511;
sine[1045] =511;
sine[1046] =511;
sine[1047] =511;
sine[1048] =511;
sine[1049] =511;
sine[1050] =511;
sine[1051] =511;
sine[1052] =511;
sine[1053] =511;
sine[1054] =511;
sine[1055] =511;
sine[1056] =511;
sine[1057] =511;
sine[1058] =511;
sine[1059] =511;
sine[1060] =511;
sine[1061] =511;
sine[1062] =511;
sine[1063] =511;
sine[1064] =511;
sine[1065] =510;
sine[1066] =510;
sine[1067] =510;
sine[1068] =510;
sine[1069] =510;
sine[1070] =510;
sine[1071] =510;
sine[1072] =510;
sine[1073] =510;
sine[1074] =510;
sine[1075] =510;
sine[1076] =510;
sine[1077] =510;
sine[1078] =510;
sine[1079] =510;
sine[1080] =510;
sine[1081] =510;
sine[1082] =510;
sine[1083] =510;
sine[1084] =510;
sine[1085] =510;
sine[1086] =510;
sine[1087] =510;
sine[1088] =510;
sine[1089] =510;
sine[1090] =510;
sine[1091] =510;
sine[1092] =510;
sine[1093] =510;
sine[1094] =510;
sine[1095] =509;
sine[1096] =509;
sine[1097] =509;
sine[1098] =509;
sine[1099] =509;
sine[1100] =509;
sine[1101] =509;
sine[1102] =509;
sine[1103] =509;
sine[1104] =509;
sine[1105] =509;
sine[1106] =509;
sine[1107] =509;
sine[1108] =509;
sine[1109] =509;
sine[1110] =509;
sine[1111] =509;
sine[1112] =509;
sine[1113] =509;
sine[1114] =509;
sine[1115] =509;
sine[1116] =508;
sine[1117] =508;
sine[1118] =508;
sine[1119] =508;
sine[1120] =508;
sine[1121] =508;
sine[1122] =508;
sine[1123] =508;
sine[1124] =508;
sine[1125] =508;
sine[1126] =508;
sine[1127] =508;
sine[1128] =508;
sine[1129] =508;
sine[1130] =508;
sine[1131] =508;
sine[1132] =508;
sine[1133] =507;
sine[1134] =507;
sine[1135] =507;
sine[1136] =507;
sine[1137] =507;
sine[1138] =507;
sine[1139] =507;
sine[1140] =507;
sine[1141] =507;
sine[1142] =507;
sine[1143] =507;
sine[1144] =507;
sine[1145] =507;
sine[1146] =507;
sine[1147] =506;
sine[1148] =506;
sine[1149] =506;
sine[1150] =506;
sine[1151] =506;
sine[1152] =506;
sine[1153] =506;
sine[1154] =506;
sine[1155] =506;
sine[1156] =506;
sine[1157] =506;
sine[1158] =506;
sine[1159] =506;
sine[1160] =505;
sine[1161] =505;
sine[1162] =505;
sine[1163] =505;
sine[1164] =505;
sine[1165] =505;
sine[1166] =505;
sine[1167] =505;
sine[1168] =505;
sine[1169] =505;
sine[1170] =505;
sine[1171] =505;
sine[1172] =504;
sine[1173] =504;
sine[1174] =504;
sine[1175] =504;
sine[1176] =504;
sine[1177] =504;
sine[1178] =504;
sine[1179] =504;
sine[1180] =504;
sine[1181] =504;
sine[1182] =504;
sine[1183] =503;
sine[1184] =503;
sine[1185] =503;
sine[1186] =503;
sine[1187] =503;
sine[1188] =503;
sine[1189] =503;
sine[1190] =503;
sine[1191] =503;
sine[1192] =503;
sine[1193] =502;
sine[1194] =502;
sine[1195] =502;
sine[1196] =502;
sine[1197] =502;
sine[1198] =502;
sine[1199] =502;
sine[1200] =502;
sine[1201] =502;
sine[1202] =502;
sine[1203] =501;
sine[1204] =501;
sine[1205] =501;
sine[1206] =501;
sine[1207] =501;
sine[1208] =501;
sine[1209] =501;
sine[1210] =501;
sine[1211] =501;
sine[1212] =500;
sine[1213] =500;
sine[1214] =500;
sine[1215] =500;
sine[1216] =500;
sine[1217] =500;
sine[1218] =500;
sine[1219] =500;
sine[1220] =500;
sine[1221] =499;
sine[1222] =499;
sine[1223] =499;
sine[1224] =499;
sine[1225] =499;
sine[1226] =499;
sine[1227] =499;
sine[1228] =499;
sine[1229] =498;
sine[1230] =498;
sine[1231] =498;
sine[1232] =498;
sine[1233] =498;
sine[1234] =498;
sine[1235] =498;
sine[1236] =498;
sine[1237] =497;
sine[1238] =497;
sine[1239] =497;
sine[1240] =497;
sine[1241] =497;
sine[1242] =497;
sine[1243] =497;
sine[1244] =497;
sine[1245] =496;
sine[1246] =496;
sine[1247] =496;
sine[1248] =496;
sine[1249] =496;
sine[1250] =496;
sine[1251] =496;
sine[1252] =496;
sine[1253] =495;
sine[1254] =495;
sine[1255] =495;
sine[1256] =495;
sine[1257] =495;
sine[1258] =495;
sine[1259] =495;
sine[1260] =494;
sine[1261] =494;
sine[1262] =494;
sine[1263] =494;
sine[1264] =494;
sine[1265] =494;
sine[1266] =494;
sine[1267] =493;
sine[1268] =493;
sine[1269] =493;
sine[1270] =493;
sine[1271] =493;
sine[1272] =493;
sine[1273] =493;
sine[1274] =492;
sine[1275] =492;
sine[1276] =492;
sine[1277] =492;
sine[1278] =492;
sine[1279] =492;
sine[1280] =492;
sine[1281] =491;
sine[1282] =491;
sine[1283] =491;
sine[1284] =491;
sine[1285] =491;
sine[1286] =491;
sine[1287] =490;
sine[1288] =490;
sine[1289] =490;
sine[1290] =490;
sine[1291] =490;
sine[1292] =490;
sine[1293] =490;
sine[1294] =489;
sine[1295] =489;
sine[1296] =489;
sine[1297] =489;
sine[1298] =489;
sine[1299] =489;
sine[1300] =488;
sine[1301] =488;
sine[1302] =488;
sine[1303] =488;
sine[1304] =488;
sine[1305] =488;
sine[1306] =487;
sine[1307] =487;
sine[1308] =487;
sine[1309] =487;
sine[1310] =487;
sine[1311] =487;
sine[1312] =486;
sine[1313] =486;
sine[1314] =486;
sine[1315] =486;
sine[1316] =486;
sine[1317] =486;
sine[1318] =485;
sine[1319] =485;
sine[1320] =485;
sine[1321] =485;
sine[1322] =485;
sine[1323] =485;
sine[1324] =484;
sine[1325] =484;
sine[1326] =484;
sine[1327] =484;
sine[1328] =484;
sine[1329] =484;
sine[1330] =483;
sine[1331] =483;
sine[1332] =483;
sine[1333] =483;
sine[1334] =483;
sine[1335] =482;
sine[1336] =482;
sine[1337] =482;
sine[1338] =482;
sine[1339] =482;
sine[1340] =482;
sine[1341] =481;
sine[1342] =481;
sine[1343] =481;
sine[1344] =481;
sine[1345] =481;
sine[1346] =480;
sine[1347] =480;
sine[1348] =480;
sine[1349] =480;
sine[1350] =480;
sine[1351] =480;
sine[1352] =479;
sine[1353] =479;
sine[1354] =479;
sine[1355] =479;
sine[1356] =479;
sine[1357] =478;
sine[1358] =478;
sine[1359] =478;
sine[1360] =478;
sine[1361] =478;
sine[1362] =477;
sine[1363] =477;
sine[1364] =477;
sine[1365] =477;
sine[1366] =477;
sine[1367] =476;
sine[1368] =476;
sine[1369] =476;
sine[1370] =476;
sine[1371] =476;
sine[1372] =475;
sine[1373] =475;
sine[1374] =475;
sine[1375] =475;
sine[1376] =475;
sine[1377] =474;
sine[1378] =474;
sine[1379] =474;
sine[1380] =474;
sine[1381] =474;
sine[1382] =473;
sine[1383] =473;
sine[1384] =473;
sine[1385] =473;
sine[1386] =473;
sine[1387] =472;
sine[1388] =472;
sine[1389] =472;
sine[1390] =472;
sine[1391] =472;
sine[1392] =471;
sine[1393] =471;
sine[1394] =471;
sine[1395] =471;
sine[1396] =471;
sine[1397] =470;
sine[1398] =470;
sine[1399] =470;
sine[1400] =470;
sine[1401] =469;
sine[1402] =469;
sine[1403] =469;
sine[1404] =469;
sine[1405] =469;
sine[1406] =468;
sine[1407] =468;
sine[1408] =468;
sine[1409] =468;
sine[1410] =468;
sine[1411] =467;
sine[1412] =467;
sine[1413] =467;
sine[1414] =467;
sine[1415] =466;
sine[1416] =466;
sine[1417] =466;
sine[1418] =466;
sine[1419] =466;
sine[1420] =465;
sine[1421] =465;
sine[1422] =465;
sine[1423] =465;
sine[1424] =464;
sine[1425] =464;
sine[1426] =464;
sine[1427] =464;
sine[1428] =463;
sine[1429] =463;
sine[1430] =463;
sine[1431] =463;
sine[1432] =463;
sine[1433] =462;
sine[1434] =462;
sine[1435] =462;
sine[1436] =462;
sine[1437] =461;
sine[1438] =461;
sine[1439] =461;
sine[1440] =461;
sine[1441] =460;
sine[1442] =460;
sine[1443] =460;
sine[1444] =460;
sine[1445] =460;
sine[1446] =459;
sine[1447] =459;
sine[1448] =459;
sine[1449] =459;
sine[1450] =458;
sine[1451] =458;
sine[1452] =458;
sine[1453] =458;
sine[1454] =457;
sine[1455] =457;
sine[1456] =457;
sine[1457] =457;
sine[1458] =456;
sine[1459] =456;
sine[1460] =456;
sine[1461] =456;
sine[1462] =455;
sine[1463] =455;
sine[1464] =455;
sine[1465] =455;
sine[1466] =454;
sine[1467] =454;
sine[1468] =454;
sine[1469] =454;
sine[1470] =454;
sine[1471] =453;
sine[1472] =453;
sine[1473] =453;
sine[1474] =453;
sine[1475] =452;
sine[1476] =452;
sine[1477] =452;
sine[1478] =452;
sine[1479] =451;
sine[1480] =451;
sine[1481] =451;
sine[1482] =450;
sine[1483] =450;
sine[1484] =450;
sine[1485] =450;
sine[1486] =449;
sine[1487] =449;
sine[1488] =449;
sine[1489] =449;
sine[1490] =448;
sine[1491] =448;
sine[1492] =448;
sine[1493] =448;
sine[1494] =447;
sine[1495] =447;
sine[1496] =447;
sine[1497] =447;
sine[1498] =446;
sine[1499] =446;
sine[1500] =446;
sine[1501] =446;
sine[1502] =445;
sine[1503] =445;
sine[1504] =445;
sine[1505] =445;
sine[1506] =444;
sine[1507] =444;
sine[1508] =444;
sine[1509] =443;
sine[1510] =443;
sine[1511] =443;
sine[1512] =443;
sine[1513] =442;
sine[1514] =442;
sine[1515] =442;
sine[1516] =442;
sine[1517] =441;
sine[1518] =441;
sine[1519] =441;
sine[1520] =441;
sine[1521] =440;
sine[1522] =440;
sine[1523] =440;
sine[1524] =439;
sine[1525] =439;
sine[1526] =439;
sine[1527] =439;
sine[1528] =438;
sine[1529] =438;
sine[1530] =438;
sine[1531] =438;
sine[1532] =437;
sine[1533] =437;
sine[1534] =437;
sine[1535] =436;
sine[1536] =436;
sine[1537] =436;
sine[1538] =436;
sine[1539] =435;
sine[1540] =435;
sine[1541] =435;
sine[1542] =434;
sine[1543] =434;
sine[1544] =434;
sine[1545] =434;
sine[1546] =433;
sine[1547] =433;
sine[1548] =433;
sine[1549] =433;
sine[1550] =432;
sine[1551] =432;
sine[1552] =432;
sine[1553] =431;
sine[1554] =431;
sine[1555] =431;
sine[1556] =431;
sine[1557] =430;
sine[1558] =430;
sine[1559] =430;
sine[1560] =429;
sine[1561] =429;
sine[1562] =429;
sine[1563] =429;
sine[1564] =428;
sine[1565] =428;
sine[1566] =428;
sine[1567] =427;
sine[1568] =427;
sine[1569] =427;
sine[1570] =427;
sine[1571] =426;
sine[1572] =426;
sine[1573] =426;
sine[1574] =425;
sine[1575] =425;
sine[1576] =425;
sine[1577] =424;
sine[1578] =424;
sine[1579] =424;
sine[1580] =424;
sine[1581] =423;
sine[1582] =423;
sine[1583] =423;
sine[1584] =422;
sine[1585] =422;
sine[1586] =422;
sine[1587] =421;
sine[1588] =421;
sine[1589] =421;
sine[1590] =421;
sine[1591] =420;
sine[1592] =420;
sine[1593] =420;
sine[1594] =419;
sine[1595] =419;
sine[1596] =419;
sine[1597] =418;
sine[1598] =418;
sine[1599] =418;
sine[1600] =418;
sine[1601] =417;
sine[1602] =417;
sine[1603] =417;
sine[1604] =416;
sine[1605] =416;
sine[1606] =416;
sine[1607] =415;
sine[1608] =415;
sine[1609] =415;
sine[1610] =415;
sine[1611] =414;
sine[1612] =414;
sine[1613] =414;
sine[1614] =413;
sine[1615] =413;
sine[1616] =413;
sine[1617] =412;
sine[1618] =412;
sine[1619] =412;
sine[1620] =411;
sine[1621] =411;
sine[1622] =411;
sine[1623] =411;
sine[1624] =410;
sine[1625] =410;
sine[1626] =410;
sine[1627] =409;
sine[1628] =409;
sine[1629] =409;
sine[1630] =408;
sine[1631] =408;
sine[1632] =408;
sine[1633] =407;
sine[1634] =407;
sine[1635] =407;
sine[1636] =406;
sine[1637] =406;
sine[1638] =406;
sine[1639] =405;
sine[1640] =405;
sine[1641] =405;
sine[1642] =405;
sine[1643] =404;
sine[1644] =404;
sine[1645] =404;
sine[1646] =403;
sine[1647] =403;
sine[1648] =403;
sine[1649] =402;
sine[1650] =402;
sine[1651] =402;
sine[1652] =401;
sine[1653] =401;
sine[1654] =401;
sine[1655] =400;
sine[1656] =400;
sine[1657] =400;
sine[1658] =399;
sine[1659] =399;
sine[1660] =399;
sine[1661] =398;
sine[1662] =398;
sine[1663] =398;
sine[1664] =397;
sine[1665] =397;
sine[1666] =397;
sine[1667] =396;
sine[1668] =396;
sine[1669] =396;
sine[1670] =395;
sine[1671] =395;
sine[1672] =395;
sine[1673] =395;
sine[1674] =394;
sine[1675] =394;
sine[1676] =394;
sine[1677] =393;
sine[1678] =393;
sine[1679] =393;
sine[1680] =392;
sine[1681] =392;
sine[1682] =392;
sine[1683] =391;
sine[1684] =391;
sine[1685] =391;
sine[1686] =390;
sine[1687] =390;
sine[1688] =390;
sine[1689] =389;
sine[1690] =389;
sine[1691] =389;
sine[1692] =388;
sine[1693] =388;
sine[1694] =388;
sine[1695] =387;
sine[1696] =387;
sine[1697] =387;
sine[1698] =386;
sine[1699] =386;
sine[1700] =386;
sine[1701] =385;
sine[1702] =385;
sine[1703] =384;
sine[1704] =384;
sine[1705] =384;
sine[1706] =383;
sine[1707] =383;
sine[1708] =383;
sine[1709] =382;
sine[1710] =382;
sine[1711] =382;
sine[1712] =381;
sine[1713] =381;
sine[1714] =381;
sine[1715] =380;
sine[1716] =380;
sine[1717] =380;
sine[1718] =379;
sine[1719] =379;
sine[1720] =379;
sine[1721] =378;
sine[1722] =378;
sine[1723] =378;
sine[1724] =377;
sine[1725] =377;
sine[1726] =377;
sine[1727] =376;
sine[1728] =376;
sine[1729] =376;
sine[1730] =375;
sine[1731] =375;
sine[1732] =375;
sine[1733] =374;
sine[1734] =374;
sine[1735] =374;
sine[1736] =373;
sine[1737] =373;
sine[1738] =372;
sine[1739] =372;
sine[1740] =372;
sine[1741] =371;
sine[1742] =371;
sine[1743] =371;
sine[1744] =370;
sine[1745] =370;
sine[1746] =370;
sine[1747] =369;
sine[1748] =369;
sine[1749] =369;
sine[1750] =368;
sine[1751] =368;
sine[1752] =368;
sine[1753] =367;
sine[1754] =367;
sine[1755] =367;
sine[1756] =366;
sine[1757] =366;
sine[1758] =365;
sine[1759] =365;
sine[1760] =365;
sine[1761] =364;
sine[1762] =364;
sine[1763] =364;
sine[1764] =363;
sine[1765] =363;
sine[1766] =363;
sine[1767] =362;
sine[1768] =362;
sine[1769] =362;
sine[1770] =361;
sine[1771] =361;
sine[1772] =360;
sine[1773] =360;
sine[1774] =360;
sine[1775] =359;
sine[1776] =359;
sine[1777] =359;
sine[1778] =358;
sine[1779] =358;
sine[1780] =358;
sine[1781] =357;
sine[1782] =357;
sine[1783] =357;
sine[1784] =356;
sine[1785] =356;
sine[1786] =355;
sine[1787] =355;
sine[1788] =355;
sine[1789] =354;
sine[1790] =354;
sine[1791] =354;
sine[1792] =353;
sine[1793] =353;
sine[1794] =353;
sine[1795] =352;
sine[1796] =352;
sine[1797] =351;
sine[1798] =351;
sine[1799] =351;
sine[1800] =350;
sine[1801] =350;
sine[1802] =350;
sine[1803] =349;
sine[1804] =349;
sine[1805] =349;
sine[1806] =348;
sine[1807] =348;
sine[1808] =347;
sine[1809] =347;
sine[1810] =347;
sine[1811] =346;
sine[1812] =346;
sine[1813] =346;
sine[1814] =345;
sine[1815] =345;
sine[1816] =345;
sine[1817] =344;
sine[1818] =344;
sine[1819] =343;
sine[1820] =343;
sine[1821] =343;
sine[1822] =342;
sine[1823] =342;
sine[1824] =342;
sine[1825] =341;
sine[1826] =341;
sine[1827] =340;
sine[1828] =340;
sine[1829] =340;
sine[1830] =339;
sine[1831] =339;
sine[1832] =339;
sine[1833] =338;
sine[1834] =338;
sine[1835] =338;
sine[1836] =337;
sine[1837] =337;
sine[1838] =336;
sine[1839] =336;
sine[1840] =336;
sine[1841] =335;
sine[1842] =335;
sine[1843] =335;
sine[1844] =334;
sine[1845] =334;
sine[1846] =333;
sine[1847] =333;
sine[1848] =333;
sine[1849] =332;
sine[1850] =332;
sine[1851] =332;
sine[1852] =331;
sine[1853] =331;
sine[1854] =330;
sine[1855] =330;
sine[1856] =330;
sine[1857] =329;
sine[1858] =329;
sine[1859] =329;
sine[1860] =328;
sine[1861] =328;
sine[1862] =327;
sine[1863] =327;
sine[1864] =327;
sine[1865] =326;
sine[1866] =326;
sine[1867] =326;
sine[1868] =325;
sine[1869] =325;
sine[1870] =324;
sine[1871] =324;
sine[1872] =324;
sine[1873] =323;
sine[1874] =323;
sine[1875] =323;
sine[1876] =322;
sine[1877] =322;
sine[1878] =321;
sine[1879] =321;
sine[1880] =321;
sine[1881] =320;
sine[1882] =320;
sine[1883] =319;
sine[1884] =319;
sine[1885] =319;
sine[1886] =318;
sine[1887] =318;
sine[1888] =318;
sine[1889] =317;
sine[1890] =317;
sine[1891] =316;
sine[1892] =316;
sine[1893] =316;
sine[1894] =315;
sine[1895] =315;
sine[1896] =315;
sine[1897] =314;
sine[1898] =314;
sine[1899] =313;
sine[1900] =313;
sine[1901] =313;
sine[1902] =312;
sine[1903] =312;
sine[1904] =311;
sine[1905] =311;
sine[1906] =311;
sine[1907] =310;
sine[1908] =310;
sine[1909] =310;
sine[1910] =309;
sine[1911] =309;
sine[1912] =308;
sine[1913] =308;
sine[1914] =308;
sine[1915] =307;
sine[1916] =307;
sine[1917] =306;
sine[1918] =306;
sine[1919] =306;
sine[1920] =305;
sine[1921] =305;
sine[1922] =305;
sine[1923] =304;
sine[1924] =304;
sine[1925] =303;
sine[1926] =303;
sine[1927] =303;
sine[1928] =302;
sine[1929] =302;
sine[1930] =301;
sine[1931] =301;
sine[1932] =301;
sine[1933] =300;
sine[1934] =300;
sine[1935] =300;
sine[1936] =299;
sine[1937] =299;
sine[1938] =298;
sine[1939] =298;
sine[1940] =298;
sine[1941] =297;
sine[1942] =297;
sine[1943] =296;
sine[1944] =296;
sine[1945] =296;
sine[1946] =295;
sine[1947] =295;
sine[1948] =295;
sine[1949] =294;
sine[1950] =294;
sine[1951] =293;
sine[1952] =293;
sine[1953] =293;
sine[1954] =292;
sine[1955] =292;
sine[1956] =291;
sine[1957] =291;
sine[1958] =291;
sine[1959] =290;
sine[1960] =290;
sine[1961] =289;
sine[1962] =289;
sine[1963] =289;
sine[1964] =288;
sine[1965] =288;
sine[1966] =288;
sine[1967] =287;
sine[1968] =287;
sine[1969] =286;
sine[1970] =286;
sine[1971] =286;
sine[1972] =285;
sine[1973] =285;
sine[1974] =284;
sine[1975] =284;
sine[1976] =284;
sine[1977] =283;
sine[1978] =283;
sine[1979] =282;
sine[1980] =282;
sine[1981] =282;
sine[1982] =281;
sine[1983] =281;
sine[1984] =281;
sine[1985] =280;
sine[1986] =280;
sine[1987] =279;
sine[1988] =279;
sine[1989] =279;
sine[1990] =278;
sine[1991] =278;
sine[1992] =277;
sine[1993] =277;
sine[1994] =277;
sine[1995] =276;
sine[1996] =276;
sine[1997] =275;
sine[1998] =275;
sine[1999] =275;
sine[2000] =274;
sine[2001] =274;
sine[2002] =274;
sine[2003] =273;
sine[2004] =273;
sine[2005] =272;
sine[2006] =272;
sine[2007] =272;
sine[2008] =271;
sine[2009] =271;
sine[2010] =270;
sine[2011] =270;
sine[2012] =270;
sine[2013] =269;
sine[2014] =269;
sine[2015] =268;
sine[2016] =268;
sine[2017] =268;
sine[2018] =267;
sine[2019] =267;
sine[2020] =266;
sine[2021] =266;
sine[2022] =266;
sine[2023] =265;
sine[2024] =265;
sine[2025] =265;
sine[2026] =264;
sine[2027] =264;
sine[2028] =263;
sine[2029] =263;
sine[2030] =263;
sine[2031] =262;
sine[2032] =262;
sine[2033] =261;
sine[2034] =261;
sine[2035] =261;
sine[2036] =260;
sine[2037] =260;
sine[2038] =259;
sine[2039] =259;
sine[2040] =259;
sine[2041] =258;
sine[2042] =258;
sine[2043] =257;
sine[2044] =257;
sine[2045] =257;
sine[2046] =256;
sine[2047] =256;
sine[2048] =256;
sine[2049] =255;
sine[2050] =255;
sine[2051] =254;
sine[2052] =254;
sine[2053] =254;
sine[2054] =253;
sine[2055] =253;
sine[2056] =252;
sine[2057] =252;
sine[2058] =252;
sine[2059] =251;
sine[2060] =251;
sine[2061] =250;
sine[2062] =250;
sine[2063] =250;
sine[2064] =249;
sine[2065] =249;
sine[2066] =248;
sine[2067] =248;
sine[2068] =248;
sine[2069] =247;
sine[2070] =247;
sine[2071] =246;
sine[2072] =246;
sine[2073] =246;
sine[2074] =245;
sine[2075] =245;
sine[2076] =245;
sine[2077] =244;
sine[2078] =244;
sine[2079] =243;
sine[2080] =243;
sine[2081] =243;
sine[2082] =242;
sine[2083] =242;
sine[2084] =241;
sine[2085] =241;
sine[2086] =241;
sine[2087] =240;
sine[2088] =240;
sine[2089] =239;
sine[2090] =239;
sine[2091] =239;
sine[2092] =238;
sine[2093] =238;
sine[2094] =237;
sine[2095] =237;
sine[2096] =237;
sine[2097] =236;
sine[2098] =236;
sine[2099] =236;
sine[2100] =235;
sine[2101] =235;
sine[2102] =234;
sine[2103] =234;
sine[2104] =234;
sine[2105] =233;
sine[2106] =233;
sine[2107] =232;
sine[2108] =232;
sine[2109] =232;
sine[2110] =231;
sine[2111] =231;
sine[2112] =230;
sine[2113] =230;
sine[2114] =230;
sine[2115] =229;
sine[2116] =229;
sine[2117] =229;
sine[2118] =228;
sine[2119] =228;
sine[2120] =227;
sine[2121] =227;
sine[2122] =227;
sine[2123] =226;
sine[2124] =226;
sine[2125] =225;
sine[2126] =225;
sine[2127] =225;
sine[2128] =224;
sine[2129] =224;
sine[2130] =223;
sine[2131] =223;
sine[2132] =223;
sine[2133] =222;
sine[2134] =222;
sine[2135] =222;
sine[2136] =221;
sine[2137] =221;
sine[2138] =220;
sine[2139] =220;
sine[2140] =220;
sine[2141] =219;
sine[2142] =219;
sine[2143] =218;
sine[2144] =218;
sine[2145] =218;
sine[2146] =217;
sine[2147] =217;
sine[2148] =216;
sine[2149] =216;
sine[2150] =216;
sine[2151] =215;
sine[2152] =215;
sine[2153] =215;
sine[2154] =214;
sine[2155] =214;
sine[2156] =213;
sine[2157] =213;
sine[2158] =213;
sine[2159] =212;
sine[2160] =212;
sine[2161] =211;
sine[2162] =211;
sine[2163] =211;
sine[2164] =210;
sine[2165] =210;
sine[2166] =210;
sine[2167] =209;
sine[2168] =209;
sine[2169] =208;
sine[2170] =208;
sine[2171] =208;
sine[2172] =207;
sine[2173] =207;
sine[2174] =206;
sine[2175] =206;
sine[2176] =206;
sine[2177] =205;
sine[2178] =205;
sine[2179] =205;
sine[2180] =204;
sine[2181] =204;
sine[2182] =203;
sine[2183] =203;
sine[2184] =203;
sine[2185] =202;
sine[2186] =202;
sine[2187] =201;
sine[2188] =201;
sine[2189] =201;
sine[2190] =200;
sine[2191] =200;
sine[2192] =200;
sine[2193] =199;
sine[2194] =199;
sine[2195] =198;
sine[2196] =198;
sine[2197] =198;
sine[2198] =197;
sine[2199] =197;
sine[2200] =196;
sine[2201] =196;
sine[2202] =196;
sine[2203] =195;
sine[2204] =195;
sine[2205] =195;
sine[2206] =194;
sine[2207] =194;
sine[2208] =193;
sine[2209] =193;
sine[2210] =193;
sine[2211] =192;
sine[2212] =192;
sine[2213] =192;
sine[2214] =191;
sine[2215] =191;
sine[2216] =190;
sine[2217] =190;
sine[2218] =190;
sine[2219] =189;
sine[2220] =189;
sine[2221] =188;
sine[2222] =188;
sine[2223] =188;
sine[2224] =187;
sine[2225] =187;
sine[2226] =187;
sine[2227] =186;
sine[2228] =186;
sine[2229] =185;
sine[2230] =185;
sine[2231] =185;
sine[2232] =184;
sine[2233] =184;
sine[2234] =184;
sine[2235] =183;
sine[2236] =183;
sine[2237] =182;
sine[2238] =182;
sine[2239] =182;
sine[2240] =181;
sine[2241] =181;
sine[2242] =181;
sine[2243] =180;
sine[2244] =180;
sine[2245] =179;
sine[2246] =179;
sine[2247] =179;
sine[2248] =178;
sine[2249] =178;
sine[2250] =178;
sine[2251] =177;
sine[2252] =177;
sine[2253] =176;
sine[2254] =176;
sine[2255] =176;
sine[2256] =175;
sine[2257] =175;
sine[2258] =175;
sine[2259] =174;
sine[2260] =174;
sine[2261] =173;
sine[2262] =173;
sine[2263] =173;
sine[2264] =172;
sine[2265] =172;
sine[2266] =172;
sine[2267] =171;
sine[2268] =171;
sine[2269] =171;
sine[2270] =170;
sine[2271] =170;
sine[2272] =169;
sine[2273] =169;
sine[2274] =169;
sine[2275] =168;
sine[2276] =168;
sine[2277] =168;
sine[2278] =167;
sine[2279] =167;
sine[2280] =166;
sine[2281] =166;
sine[2282] =166;
sine[2283] =165;
sine[2284] =165;
sine[2285] =165;
sine[2286] =164;
sine[2287] =164;
sine[2288] =164;
sine[2289] =163;
sine[2290] =163;
sine[2291] =162;
sine[2292] =162;
sine[2293] =162;
sine[2294] =161;
sine[2295] =161;
sine[2296] =161;
sine[2297] =160;
sine[2298] =160;
sine[2299] =160;
sine[2300] =159;
sine[2301] =159;
sine[2302] =158;
sine[2303] =158;
sine[2304] =158;
sine[2305] =157;
sine[2306] =157;
sine[2307] =157;
sine[2308] =156;
sine[2309] =156;
sine[2310] =156;
sine[2311] =155;
sine[2312] =155;
sine[2313] =154;
sine[2314] =154;
sine[2315] =154;
sine[2316] =153;
sine[2317] =153;
sine[2318] =153;
sine[2319] =152;
sine[2320] =152;
sine[2321] =152;
sine[2322] =151;
sine[2323] =151;
sine[2324] =151;
sine[2325] =150;
sine[2326] =150;
sine[2327] =149;
sine[2328] =149;
sine[2329] =149;
sine[2330] =148;
sine[2331] =148;
sine[2332] =148;
sine[2333] =147;
sine[2334] =147;
sine[2335] =147;
sine[2336] =146;
sine[2337] =146;
sine[2338] =146;
sine[2339] =145;
sine[2340] =145;
sine[2341] =144;
sine[2342] =144;
sine[2343] =144;
sine[2344] =143;
sine[2345] =143;
sine[2346] =143;
sine[2347] =142;
sine[2348] =142;
sine[2349] =142;
sine[2350] =141;
sine[2351] =141;
sine[2352] =141;
sine[2353] =140;
sine[2354] =140;
sine[2355] =140;
sine[2356] =139;
sine[2357] =139;
sine[2358] =139;
sine[2359] =138;
sine[2360] =138;
sine[2361] =137;
sine[2362] =137;
sine[2363] =137;
sine[2364] =136;
sine[2365] =136;
sine[2366] =136;
sine[2367] =135;
sine[2368] =135;
sine[2369] =135;
sine[2370] =134;
sine[2371] =134;
sine[2372] =134;
sine[2373] =133;
sine[2374] =133;
sine[2375] =133;
sine[2376] =132;
sine[2377] =132;
sine[2378] =132;
sine[2379] =131;
sine[2380] =131;
sine[2381] =131;
sine[2382] =130;
sine[2383] =130;
sine[2384] =130;
sine[2385] =129;
sine[2386] =129;
sine[2387] =129;
sine[2388] =128;
sine[2389] =128;
sine[2390] =128;
sine[2391] =127;
sine[2392] =127;
sine[2393] =127;
sine[2394] =126;
sine[2395] =126;
sine[2396] =125;
sine[2397] =125;
sine[2398] =125;
sine[2399] =124;
sine[2400] =124;
sine[2401] =124;
sine[2402] =123;
sine[2403] =123;
sine[2404] =123;
sine[2405] =122;
sine[2406] =122;
sine[2407] =122;
sine[2408] =121;
sine[2409] =121;
sine[2410] =121;
sine[2411] =120;
sine[2412] =120;
sine[2413] =120;
sine[2414] =119;
sine[2415] =119;
sine[2416] =119;
sine[2417] =118;
sine[2418] =118;
sine[2419] =118;
sine[2420] =117;
sine[2421] =117;
sine[2422] =117;
sine[2423] =116;
sine[2424] =116;
sine[2425] =116;
sine[2426] =116;
sine[2427] =115;
sine[2428] =115;
sine[2429] =115;
sine[2430] =114;
sine[2431] =114;
sine[2432] =114;
sine[2433] =113;
sine[2434] =113;
sine[2435] =113;
sine[2436] =112;
sine[2437] =112;
sine[2438] =112;
sine[2439] =111;
sine[2440] =111;
sine[2441] =111;
sine[2442] =110;
sine[2443] =110;
sine[2444] =110;
sine[2445] =109;
sine[2446] =109;
sine[2447] =109;
sine[2448] =108;
sine[2449] =108;
sine[2450] =108;
sine[2451] =107;
sine[2452] =107;
sine[2453] =107;
sine[2454] =106;
sine[2455] =106;
sine[2456] =106;
sine[2457] =106;
sine[2458] =105;
sine[2459] =105;
sine[2460] =105;
sine[2461] =104;
sine[2462] =104;
sine[2463] =104;
sine[2464] =103;
sine[2465] =103;
sine[2466] =103;
sine[2467] =102;
sine[2468] =102;
sine[2469] =102;
sine[2470] =101;
sine[2471] =101;
sine[2472] =101;
sine[2473] =100;
sine[2474] =100;
sine[2475] =100;
sine[2476] =100;
sine[2477] =99;
sine[2478] =99;
sine[2479] =99;
sine[2480] =98;
sine[2481] =98;
sine[2482] =98;
sine[2483] =97;
sine[2484] =97;
sine[2485] =97;
sine[2486] =96;
sine[2487] =96;
sine[2488] =96;
sine[2489] =96;
sine[2490] =95;
sine[2491] =95;
sine[2492] =95;
sine[2493] =94;
sine[2494] =94;
sine[2495] =94;
sine[2496] =93;
sine[2497] =93;
sine[2498] =93;
sine[2499] =93;
sine[2500] =92;
sine[2501] =92;
sine[2502] =92;
sine[2503] =91;
sine[2504] =91;
sine[2505] =91;
sine[2506] =90;
sine[2507] =90;
sine[2508] =90;
sine[2509] =90;
sine[2510] =89;
sine[2511] =89;
sine[2512] =89;
sine[2513] =88;
sine[2514] =88;
sine[2515] =88;
sine[2516] =87;
sine[2517] =87;
sine[2518] =87;
sine[2519] =87;
sine[2520] =86;
sine[2521] =86;
sine[2522] =86;
sine[2523] =85;
sine[2524] =85;
sine[2525] =85;
sine[2526] =84;
sine[2527] =84;
sine[2528] =84;
sine[2529] =84;
sine[2530] =83;
sine[2531] =83;
sine[2532] =83;
sine[2533] =82;
sine[2534] =82;
sine[2535] =82;
sine[2536] =82;
sine[2537] =81;
sine[2538] =81;
sine[2539] =81;
sine[2540] =80;
sine[2541] =80;
sine[2542] =80;
sine[2543] =80;
sine[2544] =79;
sine[2545] =79;
sine[2546] =79;
sine[2547] =78;
sine[2548] =78;
sine[2549] =78;
sine[2550] =78;
sine[2551] =77;
sine[2552] =77;
sine[2553] =77;
sine[2554] =77;
sine[2555] =76;
sine[2556] =76;
sine[2557] =76;
sine[2558] =75;
sine[2559] =75;
sine[2560] =75;
sine[2561] =75;
sine[2562] =74;
sine[2563] =74;
sine[2564] =74;
sine[2565] =73;
sine[2566] =73;
sine[2567] =73;
sine[2568] =73;
sine[2569] =72;
sine[2570] =72;
sine[2571] =72;
sine[2572] =72;
sine[2573] =71;
sine[2574] =71;
sine[2575] =71;
sine[2576] =70;
sine[2577] =70;
sine[2578] =70;
sine[2579] =70;
sine[2580] =69;
sine[2581] =69;
sine[2582] =69;
sine[2583] =69;
sine[2584] =68;
sine[2585] =68;
sine[2586] =68;
sine[2587] =68;
sine[2588] =67;
sine[2589] =67;
sine[2590] =67;
sine[2591] =66;
sine[2592] =66;
sine[2593] =66;
sine[2594] =66;
sine[2595] =65;
sine[2596] =65;
sine[2597] =65;
sine[2598] =65;
sine[2599] =64;
sine[2600] =64;
sine[2601] =64;
sine[2602] =64;
sine[2603] =63;
sine[2604] =63;
sine[2605] =63;
sine[2606] =63;
sine[2607] =62;
sine[2608] =62;
sine[2609] =62;
sine[2610] =62;
sine[2611] =61;
sine[2612] =61;
sine[2613] =61;
sine[2614] =61;
sine[2615] =60;
sine[2616] =60;
sine[2617] =60;
sine[2618] =59;
sine[2619] =59;
sine[2620] =59;
sine[2621] =59;
sine[2622] =58;
sine[2623] =58;
sine[2624] =58;
sine[2625] =58;
sine[2626] =57;
sine[2627] =57;
sine[2628] =57;
sine[2629] =57;
sine[2630] =57;
sine[2631] =56;
sine[2632] =56;
sine[2633] =56;
sine[2634] =56;
sine[2635] =55;
sine[2636] =55;
sine[2637] =55;
sine[2638] =55;
sine[2639] =54;
sine[2640] =54;
sine[2641] =54;
sine[2642] =54;
sine[2643] =53;
sine[2644] =53;
sine[2645] =53;
sine[2646] =53;
sine[2647] =52;
sine[2648] =52;
sine[2649] =52;
sine[2650] =52;
sine[2651] =51;
sine[2652] =51;
sine[2653] =51;
sine[2654] =51;
sine[2655] =51;
sine[2656] =50;
sine[2657] =50;
sine[2658] =50;
sine[2659] =50;
sine[2660] =49;
sine[2661] =49;
sine[2662] =49;
sine[2663] =49;
sine[2664] =48;
sine[2665] =48;
sine[2666] =48;
sine[2667] =48;
sine[2668] =48;
sine[2669] =47;
sine[2670] =47;
sine[2671] =47;
sine[2672] =47;
sine[2673] =46;
sine[2674] =46;
sine[2675] =46;
sine[2676] =46;
sine[2677] =45;
sine[2678] =45;
sine[2679] =45;
sine[2680] =45;
sine[2681] =45;
sine[2682] =44;
sine[2683] =44;
sine[2684] =44;
sine[2685] =44;
sine[2686] =43;
sine[2687] =43;
sine[2688] =43;
sine[2689] =43;
sine[2690] =43;
sine[2691] =42;
sine[2692] =42;
sine[2693] =42;
sine[2694] =42;
sine[2695] =42;
sine[2696] =41;
sine[2697] =41;
sine[2698] =41;
sine[2699] =41;
sine[2700] =40;
sine[2701] =40;
sine[2702] =40;
sine[2703] =40;
sine[2704] =40;
sine[2705] =39;
sine[2706] =39;
sine[2707] =39;
sine[2708] =39;
sine[2709] =39;
sine[2710] =38;
sine[2711] =38;
sine[2712] =38;
sine[2713] =38;
sine[2714] =38;
sine[2715] =37;
sine[2716] =37;
sine[2717] =37;
sine[2718] =37;
sine[2719] =37;
sine[2720] =36;
sine[2721] =36;
sine[2722] =36;
sine[2723] =36;
sine[2724] =36;
sine[2725] =35;
sine[2726] =35;
sine[2727] =35;
sine[2728] =35;
sine[2729] =35;
sine[2730] =34;
sine[2731] =34;
sine[2732] =34;
sine[2733] =34;
sine[2734] =34;
sine[2735] =33;
sine[2736] =33;
sine[2737] =33;
sine[2738] =33;
sine[2739] =33;
sine[2740] =32;
sine[2741] =32;
sine[2742] =32;
sine[2743] =32;
sine[2744] =32;
sine[2745] =31;
sine[2746] =31;
sine[2747] =31;
sine[2748] =31;
sine[2749] =31;
sine[2750] =31;
sine[2751] =30;
sine[2752] =30;
sine[2753] =30;
sine[2754] =30;
sine[2755] =30;
sine[2756] =29;
sine[2757] =29;
sine[2758] =29;
sine[2759] =29;
sine[2760] =29;
sine[2761] =29;
sine[2762] =28;
sine[2763] =28;
sine[2764] =28;
sine[2765] =28;
sine[2766] =28;
sine[2767] =27;
sine[2768] =27;
sine[2769] =27;
sine[2770] =27;
sine[2771] =27;
sine[2772] =27;
sine[2773] =26;
sine[2774] =26;
sine[2775] =26;
sine[2776] =26;
sine[2777] =26;
sine[2778] =26;
sine[2779] =25;
sine[2780] =25;
sine[2781] =25;
sine[2782] =25;
sine[2783] =25;
sine[2784] =25;
sine[2785] =24;
sine[2786] =24;
sine[2787] =24;
sine[2788] =24;
sine[2789] =24;
sine[2790] =24;
sine[2791] =23;
sine[2792] =23;
sine[2793] =23;
sine[2794] =23;
sine[2795] =23;
sine[2796] =23;
sine[2797] =22;
sine[2798] =22;
sine[2799] =22;
sine[2800] =22;
sine[2801] =22;
sine[2802] =22;
sine[2803] =21;
sine[2804] =21;
sine[2805] =21;
sine[2806] =21;
sine[2807] =21;
sine[2808] =21;
sine[2809] =21;
sine[2810] =20;
sine[2811] =20;
sine[2812] =20;
sine[2813] =20;
sine[2814] =20;
sine[2815] =20;
sine[2816] =19;
sine[2817] =19;
sine[2818] =19;
sine[2819] =19;
sine[2820] =19;
sine[2821] =19;
sine[2822] =19;
sine[2823] =18;
sine[2824] =18;
sine[2825] =18;
sine[2826] =18;
sine[2827] =18;
sine[2828] =18;
sine[2829] =18;
sine[2830] =17;
sine[2831] =17;
sine[2832] =17;
sine[2833] =17;
sine[2834] =17;
sine[2835] =17;
sine[2836] =17;
sine[2837] =16;
sine[2838] =16;
sine[2839] =16;
sine[2840] =16;
sine[2841] =16;
sine[2842] =16;
sine[2843] =16;
sine[2844] =15;
sine[2845] =15;
sine[2846] =15;
sine[2847] =15;
sine[2848] =15;
sine[2849] =15;
sine[2850] =15;
sine[2851] =15;
sine[2852] =14;
sine[2853] =14;
sine[2854] =14;
sine[2855] =14;
sine[2856] =14;
sine[2857] =14;
sine[2858] =14;
sine[2859] =14;
sine[2860] =13;
sine[2861] =13;
sine[2862] =13;
sine[2863] =13;
sine[2864] =13;
sine[2865] =13;
sine[2866] =13;
sine[2867] =13;
sine[2868] =12;
sine[2869] =12;
sine[2870] =12;
sine[2871] =12;
sine[2872] =12;
sine[2873] =12;
sine[2874] =12;
sine[2875] =12;
sine[2876] =11;
sine[2877] =11;
sine[2878] =11;
sine[2879] =11;
sine[2880] =11;
sine[2881] =11;
sine[2882] =11;
sine[2883] =11;
sine[2884] =11;
sine[2885] =10;
sine[2886] =10;
sine[2887] =10;
sine[2888] =10;
sine[2889] =10;
sine[2890] =10;
sine[2891] =10;
sine[2892] =10;
sine[2893] =10;
sine[2894] =9;
sine[2895] =9;
sine[2896] =9;
sine[2897] =9;
sine[2898] =9;
sine[2899] =9;
sine[2900] =9;
sine[2901] =9;
sine[2902] =9;
sine[2903] =9;
sine[2904] =8;
sine[2905] =8;
sine[2906] =8;
sine[2907] =8;
sine[2908] =8;
sine[2909] =8;
sine[2910] =8;
sine[2911] =8;
sine[2912] =8;
sine[2913] =8;
sine[2914] =7;
sine[2915] =7;
sine[2916] =7;
sine[2917] =7;
sine[2918] =7;
sine[2919] =7;
sine[2920] =7;
sine[2921] =7;
sine[2922] =7;
sine[2923] =7;
sine[2924] =7;
sine[2925] =6;
sine[2926] =6;
sine[2927] =6;
sine[2928] =6;
sine[2929] =6;
sine[2930] =6;
sine[2931] =6;
sine[2932] =6;
sine[2933] =6;
sine[2934] =6;
sine[2935] =6;
sine[2936] =6;
sine[2937] =5;
sine[2938] =5;
sine[2939] =5;
sine[2940] =5;
sine[2941] =5;
sine[2942] =5;
sine[2943] =5;
sine[2944] =5;
sine[2945] =5;
sine[2946] =5;
sine[2947] =5;
sine[2948] =5;
sine[2949] =5;
sine[2950] =4;
sine[2951] =4;
sine[2952] =4;
sine[2953] =4;
sine[2954] =4;
sine[2955] =4;
sine[2956] =4;
sine[2957] =4;
sine[2958] =4;
sine[2959] =4;
sine[2960] =4;
sine[2961] =4;
sine[2962] =4;
sine[2963] =4;
sine[2964] =3;
sine[2965] =3;
sine[2966] =3;
sine[2967] =3;
sine[2968] =3;
sine[2969] =3;
sine[2970] =3;
sine[2971] =3;
sine[2972] =3;
sine[2973] =3;
sine[2974] =3;
sine[2975] =3;
sine[2976] =3;
sine[2977] =3;
sine[2978] =3;
sine[2979] =3;
sine[2980] =3;
sine[2981] =2;
sine[2982] =2;
sine[2983] =2;
sine[2984] =2;
sine[2985] =2;
sine[2986] =2;
sine[2987] =2;
sine[2988] =2;
sine[2989] =2;
sine[2990] =2;
sine[2991] =2;
sine[2992] =2;
sine[2993] =2;
sine[2994] =2;
sine[2995] =2;
sine[2996] =2;
sine[2997] =2;
sine[2998] =2;
sine[2999] =2;
sine[3000] =2;
sine[3001] =2;
sine[3002] =1;
sine[3003] =1;
sine[3004] =1;
sine[3005] =1;
sine[3006] =1;
sine[3007] =1;
sine[3008] =1;
sine[3009] =1;
sine[3010] =1;
sine[3011] =1;
sine[3012] =1;
sine[3013] =1;
sine[3014] =1;
sine[3015] =1;
sine[3016] =1;
sine[3017] =1;
sine[3018] =1;
sine[3019] =1;
sine[3020] =1;
sine[3021] =1;
sine[3022] =1;
sine[3023] =1;
sine[3024] =1;
sine[3025] =1;
sine[3026] =1;
sine[3027] =1;
sine[3028] =1;
sine[3029] =1;
sine[3030] =1;
sine[3031] =1;
sine[3032] =0;
sine[3033] =0;
sine[3034] =0;
sine[3035] =0;
sine[3036] =0;
sine[3037] =0;
sine[3038] =0;
sine[3039] =0;
sine[3040] =0;
sine[3041] =0;
sine[3042] =0;
sine[3043] =0;
sine[3044] =0;
sine[3045] =0;
sine[3046] =0;
sine[3047] =0;
sine[3048] =0;
sine[3049] =0;
sine[3050] =0;
sine[3051] =0;
sine[3052] =0;
sine[3053] =0;
sine[3054] =0;
sine[3055] =0;
sine[3056] =0;
sine[3057] =0;
sine[3058] =0;
sine[3059] =0;
sine[3060] =0;
sine[3061] =0;
sine[3062] =0;
sine[3063] =0;
sine[3064] =0;
sine[3065] =0;
sine[3066] =0;
sine[3067] =0;
sine[3068] =0;
sine[3069] =0;
sine[3070] =0;
sine[3071] =0;
sine[3072] =0;
sine[3073] =0;
sine[3074] =0;
sine[3075] =0;
sine[3076] =0;
sine[3077] =0;
sine[3078] =0;
sine[3079] =0;
sine[3080] =0;
sine[3081] =0;
sine[3082] =0;
sine[3083] =0;
sine[3084] =0;
sine[3085] =0;
sine[3086] =0;
sine[3087] =0;
sine[3088] =0;
sine[3089] =0;
sine[3090] =0;
sine[3091] =0;
sine[3092] =0;
sine[3093] =0;
sine[3094] =0;
sine[3095] =0;
sine[3096] =0;
sine[3097] =0;
sine[3098] =0;
sine[3099] =0;
sine[3100] =0;
sine[3101] =0;
sine[3102] =0;
sine[3103] =0;
sine[3104] =0;
sine[3105] =0;
sine[3106] =0;
sine[3107] =0;
sine[3108] =0;
sine[3109] =0;
sine[3110] =0;
sine[3111] =0;
sine[3112] =0;
sine[3113] =1;
sine[3114] =1;
sine[3115] =1;
sine[3116] =1;
sine[3117] =1;
sine[3118] =1;
sine[3119] =1;
sine[3120] =1;
sine[3121] =1;
sine[3122] =1;
sine[3123] =1;
sine[3124] =1;
sine[3125] =1;
sine[3126] =1;
sine[3127] =1;
sine[3128] =1;
sine[3129] =1;
sine[3130] =1;
sine[3131] =1;
sine[3132] =1;
sine[3133] =1;
sine[3134] =1;
sine[3135] =1;
sine[3136] =1;
sine[3137] =1;
sine[3138] =1;
sine[3139] =1;
sine[3140] =1;
sine[3141] =1;
sine[3142] =1;
sine[3143] =2;
sine[3144] =2;
sine[3145] =2;
sine[3146] =2;
sine[3147] =2;
sine[3148] =2;
sine[3149] =2;
sine[3150] =2;
sine[3151] =2;
sine[3152] =2;
sine[3153] =2;
sine[3154] =2;
sine[3155] =2;
sine[3156] =2;
sine[3157] =2;
sine[3158] =2;
sine[3159] =2;
sine[3160] =2;
sine[3161] =2;
sine[3162] =2;
sine[3163] =2;
sine[3164] =3;
sine[3165] =3;
sine[3166] =3;
sine[3167] =3;
sine[3168] =3;
sine[3169] =3;
sine[3170] =3;
sine[3171] =3;
sine[3172] =3;
sine[3173] =3;
sine[3174] =3;
sine[3175] =3;
sine[3176] =3;
sine[3177] =3;
sine[3178] =3;
sine[3179] =3;
sine[3180] =3;
sine[3181] =4;
sine[3182] =4;
sine[3183] =4;
sine[3184] =4;
sine[3185] =4;
sine[3186] =4;
sine[3187] =4;
sine[3188] =4;
sine[3189] =4;
sine[3190] =4;
sine[3191] =4;
sine[3192] =4;
sine[3193] =4;
sine[3194] =4;
sine[3195] =5;
sine[3196] =5;
sine[3197] =5;
sine[3198] =5;
sine[3199] =5;
sine[3200] =5;
sine[3201] =5;
sine[3202] =5;
sine[3203] =5;
sine[3204] =5;
sine[3205] =5;
sine[3206] =5;
sine[3207] =5;
sine[3208] =6;
sine[3209] =6;
sine[3210] =6;
sine[3211] =6;
sine[3212] =6;
sine[3213] =6;
sine[3214] =6;
sine[3215] =6;
sine[3216] =6;
sine[3217] =6;
sine[3218] =6;
sine[3219] =6;
sine[3220] =7;
sine[3221] =7;
sine[3222] =7;
sine[3223] =7;
sine[3224] =7;
sine[3225] =7;
sine[3226] =7;
sine[3227] =7;
sine[3228] =7;
sine[3229] =7;
sine[3230] =7;
sine[3231] =8;
sine[3232] =8;
sine[3233] =8;
sine[3234] =8;
sine[3235] =8;
sine[3236] =8;
sine[3237] =8;
sine[3238] =8;
sine[3239] =8;
sine[3240] =8;
sine[3241] =9;
sine[3242] =9;
sine[3243] =9;
sine[3244] =9;
sine[3245] =9;
sine[3246] =9;
sine[3247] =9;
sine[3248] =9;
sine[3249] =9;
sine[3250] =9;
sine[3251] =10;
sine[3252] =10;
sine[3253] =10;
sine[3254] =10;
sine[3255] =10;
sine[3256] =10;
sine[3257] =10;
sine[3258] =10;
sine[3259] =10;
sine[3260] =11;
sine[3261] =11;
sine[3262] =11;
sine[3263] =11;
sine[3264] =11;
sine[3265] =11;
sine[3266] =11;
sine[3267] =11;
sine[3268] =11;
sine[3269] =12;
sine[3270] =12;
sine[3271] =12;
sine[3272] =12;
sine[3273] =12;
sine[3274] =12;
sine[3275] =12;
sine[3276] =12;
sine[3277] =13;
sine[3278] =13;
sine[3279] =13;
sine[3280] =13;
sine[3281] =13;
sine[3282] =13;
sine[3283] =13;
sine[3284] =13;
sine[3285] =14;
sine[3286] =14;
sine[3287] =14;
sine[3288] =14;
sine[3289] =14;
sine[3290] =14;
sine[3291] =14;
sine[3292] =14;
sine[3293] =15;
sine[3294] =15;
sine[3295] =15;
sine[3296] =15;
sine[3297] =15;
sine[3298] =15;
sine[3299] =15;
sine[3300] =15;
sine[3301] =16;
sine[3302] =16;
sine[3303] =16;
sine[3304] =16;
sine[3305] =16;
sine[3306] =16;
sine[3307] =16;
sine[3308] =17;
sine[3309] =17;
sine[3310] =17;
sine[3311] =17;
sine[3312] =17;
sine[3313] =17;
sine[3314] =17;
sine[3315] =18;
sine[3316] =18;
sine[3317] =18;
sine[3318] =18;
sine[3319] =18;
sine[3320] =18;
sine[3321] =18;
sine[3322] =19;
sine[3323] =19;
sine[3324] =19;
sine[3325] =19;
sine[3326] =19;
sine[3327] =19;
sine[3328] =19;
sine[3329] =20;
sine[3330] =20;
sine[3331] =20;
sine[3332] =20;
sine[3333] =20;
sine[3334] =20;
sine[3335] =21;
sine[3336] =21;
sine[3337] =21;
sine[3338] =21;
sine[3339] =21;
sine[3340] =21;
sine[3341] =21;
sine[3342] =22;
sine[3343] =22;
sine[3344] =22;
sine[3345] =22;
sine[3346] =22;
sine[3347] =22;
sine[3348] =23;
sine[3349] =23;
sine[3350] =23;
sine[3351] =23;
sine[3352] =23;
sine[3353] =23;
sine[3354] =24;
sine[3355] =24;
sine[3356] =24;
sine[3357] =24;
sine[3358] =24;
sine[3359] =24;
sine[3360] =25;
sine[3361] =25;
sine[3362] =25;
sine[3363] =25;
sine[3364] =25;
sine[3365] =25;
sine[3366] =26;
sine[3367] =26;
sine[3368] =26;
sine[3369] =26;
sine[3370] =26;
sine[3371] =26;
sine[3372] =27;
sine[3373] =27;
sine[3374] =27;
sine[3375] =27;
sine[3376] =27;
sine[3377] =27;
sine[3378] =28;
sine[3379] =28;
sine[3380] =28;
sine[3381] =28;
sine[3382] =28;
sine[3383] =29;
sine[3384] =29;
sine[3385] =29;
sine[3386] =29;
sine[3387] =29;
sine[3388] =29;
sine[3389] =30;
sine[3390] =30;
sine[3391] =30;
sine[3392] =30;
sine[3393] =30;
sine[3394] =31;
sine[3395] =31;
sine[3396] =31;
sine[3397] =31;
sine[3398] =31;
sine[3399] =31;
sine[3400] =32;
sine[3401] =32;
sine[3402] =32;
sine[3403] =32;
sine[3404] =32;
sine[3405] =33;
sine[3406] =33;
sine[3407] =33;
sine[3408] =33;
sine[3409] =33;
sine[3410] =34;
sine[3411] =34;
sine[3412] =34;
sine[3413] =34;
sine[3414] =34;
sine[3415] =35;
sine[3416] =35;
sine[3417] =35;
sine[3418] =35;
sine[3419] =35;
sine[3420] =36;
sine[3421] =36;
sine[3422] =36;
sine[3423] =36;
sine[3424] =36;
sine[3425] =37;
sine[3426] =37;
sine[3427] =37;
sine[3428] =37;
sine[3429] =37;
sine[3430] =38;
sine[3431] =38;
sine[3432] =38;
sine[3433] =38;
sine[3434] =38;
sine[3435] =39;
sine[3436] =39;
sine[3437] =39;
sine[3438] =39;
sine[3439] =39;
sine[3440] =40;
sine[3441] =40;
sine[3442] =40;
sine[3443] =40;
sine[3444] =40;
sine[3445] =41;
sine[3446] =41;
sine[3447] =41;
sine[3448] =41;
sine[3449] =42;
sine[3450] =42;
sine[3451] =42;
sine[3452] =42;
sine[3453] =42;
sine[3454] =43;
sine[3455] =43;
sine[3456] =43;
sine[3457] =43;
sine[3458] =43;
sine[3459] =44;
sine[3460] =44;
sine[3461] =44;
sine[3462] =44;
sine[3463] =45;
sine[3464] =45;
sine[3465] =45;
sine[3466] =45;
sine[3467] =45;
sine[3468] =46;
sine[3469] =46;
sine[3470] =46;
sine[3471] =46;
sine[3472] =47;
sine[3473] =47;
sine[3474] =47;
sine[3475] =47;
sine[3476] =48;
sine[3477] =48;
sine[3478] =48;
sine[3479] =48;
sine[3480] =48;
sine[3481] =49;
sine[3482] =49;
sine[3483] =49;
sine[3484] =49;
sine[3485] =50;
sine[3486] =50;
sine[3487] =50;
sine[3488] =50;
sine[3489] =51;
sine[3490] =51;
sine[3491] =51;
sine[3492] =51;
sine[3493] =51;
sine[3494] =52;
sine[3495] =52;
sine[3496] =52;
sine[3497] =52;
sine[3498] =53;
sine[3499] =53;
sine[3500] =53;
sine[3501] =53;
sine[3502] =54;
sine[3503] =54;
sine[3504] =54;
sine[3505] =54;
sine[3506] =55;
sine[3507] =55;
sine[3508] =55;
sine[3509] =55;
sine[3510] =56;
sine[3511] =56;
sine[3512] =56;
sine[3513] =56;
sine[3514] =57;
sine[3515] =57;
sine[3516] =57;
sine[3517] =57;
sine[3518] =57;
sine[3519] =58;
sine[3520] =58;
sine[3521] =58;
sine[3522] =58;
sine[3523] =59;
sine[3524] =59;
sine[3525] =59;
sine[3526] =59;
sine[3527] =60;
sine[3528] =60;
sine[3529] =60;
sine[3530] =61;
sine[3531] =61;
sine[3532] =61;
sine[3533] =61;
sine[3534] =62;
sine[3535] =62;
sine[3536] =62;
sine[3537] =62;
sine[3538] =63;
sine[3539] =63;
sine[3540] =63;
sine[3541] =63;
sine[3542] =64;
sine[3543] =64;
sine[3544] =64;
sine[3545] =64;
sine[3546] =65;
sine[3547] =65;
sine[3548] =65;
sine[3549] =65;
sine[3550] =66;
sine[3551] =66;
sine[3552] =66;
sine[3553] =66;
sine[3554] =67;
sine[3555] =67;
sine[3556] =67;
sine[3557] =68;
sine[3558] =68;
sine[3559] =68;
sine[3560] =68;
sine[3561] =69;
sine[3562] =69;
sine[3563] =69;
sine[3564] =69;
sine[3565] =70;
sine[3566] =70;
sine[3567] =70;
sine[3568] =70;
sine[3569] =71;
sine[3570] =71;
sine[3571] =71;
sine[3572] =72;
sine[3573] =72;
sine[3574] =72;
sine[3575] =72;
sine[3576] =73;
sine[3577] =73;
sine[3578] =73;
sine[3579] =73;
sine[3580] =74;
sine[3581] =74;
sine[3582] =74;
sine[3583] =75;
sine[3584] =75;
sine[3585] =75;
sine[3586] =75;
sine[3587] =76;
sine[3588] =76;
sine[3589] =76;
sine[3590] =77;
sine[3591] =77;
sine[3592] =77;
sine[3593] =77;
sine[3594] =78;
sine[3595] =78;
sine[3596] =78;
sine[3597] =78;
sine[3598] =79;
sine[3599] =79;
sine[3600] =79;
sine[3601] =80;
sine[3602] =80;
sine[3603] =80;
sine[3604] =80;
sine[3605] =81;
sine[3606] =81;
sine[3607] =81;
sine[3608] =82;
sine[3609] =82;
sine[3610] =82;
sine[3611] =82;
sine[3612] =83;
sine[3613] =83;
sine[3614] =83;
sine[3615] =84;
sine[3616] =84;
sine[3617] =84;
sine[3618] =84;
sine[3619] =85;
sine[3620] =85;
sine[3621] =85;
sine[3622] =86;
sine[3623] =86;
sine[3624] =86;
sine[3625] =87;
sine[3626] =87;
sine[3627] =87;
sine[3628] =87;
sine[3629] =88;
sine[3630] =88;
sine[3631] =88;
sine[3632] =89;
sine[3633] =89;
sine[3634] =89;
sine[3635] =90;
sine[3636] =90;
sine[3637] =90;
sine[3638] =90;
sine[3639] =91;
sine[3640] =91;
sine[3641] =91;
sine[3642] =92;
sine[3643] =92;
sine[3644] =92;
sine[3645] =93;
sine[3646] =93;
sine[3647] =93;
sine[3648] =93;
sine[3649] =94;
sine[3650] =94;
sine[3651] =94;
sine[3652] =95;
sine[3653] =95;
sine[3654] =95;
sine[3655] =96;
sine[3656] =96;
sine[3657] =96;
sine[3658] =96;
sine[3659] =97;
sine[3660] =97;
sine[3661] =97;
sine[3662] =98;
sine[3663] =98;
sine[3664] =98;
sine[3665] =99;
sine[3666] =99;
sine[3667] =99;
sine[3668] =100;
sine[3669] =100;
sine[3670] =100;
sine[3671] =100;
sine[3672] =101;
sine[3673] =101;
sine[3674] =101;
sine[3675] =102;
sine[3676] =102;
sine[3677] =102;
sine[3678] =103;
sine[3679] =103;
sine[3680] =103;
sine[3681] =104;
sine[3682] =104;
sine[3683] =104;
sine[3684] =105;
sine[3685] =105;
sine[3686] =105;
sine[3687] =106;
sine[3688] =106;
sine[3689] =106;
sine[3690] =106;
sine[3691] =107;
sine[3692] =107;
sine[3693] =107;
sine[3694] =108;
sine[3695] =108;
sine[3696] =108;
sine[3697] =109;
sine[3698] =109;
sine[3699] =109;
sine[3700] =110;
sine[3701] =110;
sine[3702] =110;
sine[3703] =111;
sine[3704] =111;
sine[3705] =111;
sine[3706] =112;
sine[3707] =112;
sine[3708] =112;
sine[3709] =113;
sine[3710] =113;
sine[3711] =113;
sine[3712] =114;
sine[3713] =114;
sine[3714] =114;
sine[3715] =115;
sine[3716] =115;
sine[3717] =115;
sine[3718] =116;
sine[3719] =116;
sine[3720] =116;
sine[3721] =116;
sine[3722] =117;
sine[3723] =117;
sine[3724] =117;
sine[3725] =118;
sine[3726] =118;
sine[3727] =118;
sine[3728] =119;
sine[3729] =119;
sine[3730] =119;
sine[3731] =120;
sine[3732] =120;
sine[3733] =120;
sine[3734] =121;
sine[3735] =121;
sine[3736] =121;
sine[3737] =122;
sine[3738] =122;
sine[3739] =122;
sine[3740] =123;
sine[3741] =123;
sine[3742] =123;
sine[3743] =124;
sine[3744] =124;
sine[3745] =124;
sine[3746] =125;
sine[3747] =125;
sine[3748] =125;
sine[3749] =126;
sine[3750] =126;
sine[3751] =127;
sine[3752] =127;
sine[3753] =127;
sine[3754] =128;
sine[3755] =128;
sine[3756] =128;
sine[3757] =129;
sine[3758] =129;
sine[3759] =129;
sine[3760] =130;
sine[3761] =130;
sine[3762] =130;
sine[3763] =131;
sine[3764] =131;
sine[3765] =131;
sine[3766] =132;
sine[3767] =132;
sine[3768] =132;
sine[3769] =133;
sine[3770] =133;
sine[3771] =133;
sine[3772] =134;
sine[3773] =134;
sine[3774] =134;
sine[3775] =135;
sine[3776] =135;
sine[3777] =135;
sine[3778] =136;
sine[3779] =136;
sine[3780] =136;
sine[3781] =137;
sine[3782] =137;
sine[3783] =137;
sine[3784] =138;
sine[3785] =138;
sine[3786] =139;
sine[3787] =139;
sine[3788] =139;
sine[3789] =140;
sine[3790] =140;
sine[3791] =140;
sine[3792] =141;
sine[3793] =141;
sine[3794] =141;
sine[3795] =142;
sine[3796] =142;
sine[3797] =142;
sine[3798] =143;
sine[3799] =143;
sine[3800] =143;
sine[3801] =144;
sine[3802] =144;
sine[3803] =144;
sine[3804] =145;
sine[3805] =145;
sine[3806] =146;
sine[3807] =146;
sine[3808] =146;
sine[3809] =147;
sine[3810] =147;
sine[3811] =147;
sine[3812] =148;
sine[3813] =148;
sine[3814] =148;
sine[3815] =149;
sine[3816] =149;
sine[3817] =149;
sine[3818] =150;
sine[3819] =150;
sine[3820] =151;
sine[3821] =151;
sine[3822] =151;
sine[3823] =152;
sine[3824] =152;
sine[3825] =152;
sine[3826] =153;
sine[3827] =153;
sine[3828] =153;
sine[3829] =154;
sine[3830] =154;
sine[3831] =154;
sine[3832] =155;
sine[3833] =155;
sine[3834] =156;
sine[3835] =156;
sine[3836] =156;
sine[3837] =157;
sine[3838] =157;
sine[3839] =157;
sine[3840] =158;
sine[3841] =158;
sine[3842] =158;
sine[3843] =159;
sine[3844] =159;
sine[3845] =160;
sine[3846] =160;
sine[3847] =160;
sine[3848] =161;
sine[3849] =161;
sine[3850] =161;
sine[3851] =162;
sine[3852] =162;
sine[3853] =162;
sine[3854] =163;
sine[3855] =163;
sine[3856] =164;
sine[3857] =164;
sine[3858] =164;
sine[3859] =165;
sine[3860] =165;
sine[3861] =165;
sine[3862] =166;
sine[3863] =166;
sine[3864] =166;
sine[3865] =167;
sine[3866] =167;
sine[3867] =168;
sine[3868] =168;
sine[3869] =168;
sine[3870] =169;
sine[3871] =169;
sine[3872] =169;
sine[3873] =170;
sine[3874] =170;
sine[3875] =171;
sine[3876] =171;
sine[3877] =171;
sine[3878] =172;
sine[3879] =172;
sine[3880] =172;
sine[3881] =173;
sine[3882] =173;
sine[3883] =173;
sine[3884] =174;
sine[3885] =174;
sine[3886] =175;
sine[3887] =175;
sine[3888] =175;
sine[3889] =176;
sine[3890] =176;
sine[3891] =176;
sine[3892] =177;
sine[3893] =177;
sine[3894] =178;
sine[3895] =178;
sine[3896] =178;
sine[3897] =179;
sine[3898] =179;
sine[3899] =179;
sine[3900] =180;
sine[3901] =180;
sine[3902] =181;
sine[3903] =181;
sine[3904] =181;
sine[3905] =182;
sine[3906] =182;
sine[3907] =182;
sine[3908] =183;
sine[3909] =183;
sine[3910] =184;
sine[3911] =184;
sine[3912] =184;
sine[3913] =185;
sine[3914] =185;
sine[3915] =185;
sine[3916] =186;
sine[3917] =186;
sine[3918] =187;
sine[3919] =187;
sine[3920] =187;
sine[3921] =188;
sine[3922] =188;
sine[3923] =188;
sine[3924] =189;
sine[3925] =189;
sine[3926] =190;
sine[3927] =190;
sine[3928] =190;
sine[3929] =191;
sine[3930] =191;
sine[3931] =192;
sine[3932] =192;
sine[3933] =192;
sine[3934] =193;
sine[3935] =193;
sine[3936] =193;
sine[3937] =194;
sine[3938] =194;
sine[3939] =195;
sine[3940] =195;
sine[3941] =195;
sine[3942] =196;
sine[3943] =196;
sine[3944] =196;
sine[3945] =197;
sine[3946] =197;
sine[3947] =198;
sine[3948] =198;
sine[3949] =198;
sine[3950] =199;
sine[3951] =199;
sine[3952] =200;
sine[3953] =200;
sine[3954] =200;
sine[3955] =201;
sine[3956] =201;
sine[3957] =201;
sine[3958] =202;
sine[3959] =202;
sine[3960] =203;
sine[3961] =203;
sine[3962] =203;
sine[3963] =204;
sine[3964] =204;
sine[3965] =205;
sine[3966] =205;
sine[3967] =205;
sine[3968] =206;
sine[3969] =206;
sine[3970] =206;
sine[3971] =207;
sine[3972] =207;
sine[3973] =208;
sine[3974] =208;
sine[3975] =208;
sine[3976] =209;
sine[3977] =209;
sine[3978] =210;
sine[3979] =210;
sine[3980] =210;
sine[3981] =211;
sine[3982] =211;
sine[3983] =211;
sine[3984] =212;
sine[3985] =212;
sine[3986] =213;
sine[3987] =213;
sine[3988] =213;
sine[3989] =214;
sine[3990] =214;
sine[3991] =215;
sine[3992] =215;
sine[3993] =215;
sine[3994] =216;
sine[3995] =216;
sine[3996] =216;
sine[3997] =217;
sine[3998] =217;
sine[3999] =218;
sine[4000] =218;
sine[4001] =218;
sine[4002] =219;
sine[4003] =219;
sine[4004] =220;
sine[4005] =220;
sine[4006] =220;
sine[4007] =221;
sine[4008] =221;
sine[4009] =222;
sine[4010] =222;
sine[4011] =222;
sine[4012] =223;
sine[4013] =223;
sine[4014] =223;
sine[4015] =224;
sine[4016] =224;
sine[4017] =225;
sine[4018] =225;
sine[4019] =225;
sine[4020] =226;
sine[4021] =226;
sine[4022] =227;
sine[4023] =227;
sine[4024] =227;
sine[4025] =228;
sine[4026] =228;
sine[4027] =229;
sine[4028] =229;
sine[4029] =229;
sine[4030] =230;
sine[4031] =230;
sine[4032] =230;
sine[4033] =231;
sine[4034] =231;
sine[4035] =232;
sine[4036] =232;
sine[4037] =232;
sine[4038] =233;
sine[4039] =233;
sine[4040] =234;
sine[4041] =234;
sine[4042] =234;
sine[4043] =235;
sine[4044] =235;
sine[4045] =236;
sine[4046] =236;
sine[4047] =236;
sine[4048] =237;
sine[4049] =237;
sine[4050] =237;
sine[4051] =238;
sine[4052] =238;
sine[4053] =239;
sine[4054] =239;
sine[4055] =239;
sine[4056] =240;
sine[4057] =240;
sine[4058] =241;
sine[4059] =241;
sine[4060] =241;
sine[4061] =242;
sine[4062] =242;
sine[4063] =243;
sine[4064] =243;
sine[4065] =243;
sine[4066] =244;
sine[4067] =244;
sine[4068] =245;
sine[4069] =245;
sine[4070] =245;
sine[4071] =246;
sine[4072] =246;
sine[4073] =246;
sine[4074] =247;
sine[4075] =247;
sine[4076] =248;
sine[4077] =248;
sine[4078] =248;
sine[4079] =249;
sine[4080] =249;
sine[4081] =250;
sine[4082] =250;
sine[4083] =250;
sine[4084] =251;
sine[4085] =251;
sine[4086] =252;
sine[4087] =252;
sine[4088] =252;
sine[4089] =253;
sine[4090] =253;
sine[4091] =254;
sine[4092] =254;
sine[4093] =254;
sine[4094] =255;
sine[4095] =255;

    end
    always@ (posedge(Clk))
    begin
        data_out_1 = sine[i];
        i = i+ 1;
        if(i == 4095)
            i = 0;
    end
endmodule